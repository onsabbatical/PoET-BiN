--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:24:12 07/23/2019
-- Design Name:   
-- Module Name:   D:/siva/Masters/Thesis/07_ETE_19/part_svhn/cifar_rinc_40_8_tb.vhd
-- Project Name:  part_svhn
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: cifar_rinc_40_8
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY cifar_rinc_40_8_tb IS
END cifar_rinc_40_8_tb;
 
ARCHITECTURE behavior OF cifar_rinc_40_8_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT cifar_rinc_40_8
    PORT(
         inp_feat : IN  std_logic_vector(511 downto 0);
			cor_out :OUT std_logic_vector(79 downto 0);
			cor_in : IN std_logic_vector(79 downto 0);
         pred_out : OUT  std_logic_vector(79 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal inp_feat : std_logic_vector(511 downto 0) := (others => '0');
	signal cor_in : std_logic_vector(79 downto 0) := (others => '0');

 	--Outputs
   signal pred_out : std_logic_vector(79 downto 0);
	signal cor_out : std_logic_vector(79 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   -- constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: cifar_rinc_40_8 PORT MAP (
          inp_feat => inp_feat,
			 cor_out => cor_out,
			 cor_in => cor_in,
          pred_out => pred_out
        );

   -- Clock process definitions
   -- <clock>_process :process
   -- begin
		-- <clock> <= '0';
		-- wait for <clock>_period/2;
		-- <clock> <= '1';
		-- wait for <clock>_period/2;
   -- end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      -- wait for <clock>_period*10;
inp_feat <= "11111111111111110011010110011111111111110001011011101010011110110111111111111001111111111111111101100111111111011111011111100111111111011111111111111110111111111011100111100011011111010101011111110110011111010010010010110100111111100101111111111011111111111000100111110001101101011000110101010111111100011111111111111111111110011110101111100101100111110100101101111101111101111110100011100101011011111010001101110101010111011101110111110110111011111111111010111111101111010101101111011000100010010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110111011111011110110010110111111111111111111111011111010101111011110111110101011101111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111111111010110111101101101110011110011011111111111111001010110111101110111100111010111101101111111001101011011111101011110001111111101111111011110111111101111010101111111011111011111101111111101111111111111111010001111101111111001110111101101110001111011100111101110110110101111111110110101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011111110011111011111111010100111111111111110011111111111011101111011111111110101011101111101111010111111111110101101111111110011111111101111111011000010111010000101011111001111111111010110111101101111110110110011111111111111111001011110111101110111111111010111101101111111001100011011111101011110001011011101111111011110111111001101011101111111011111111111101111111101111111111111111010101111101111110001110111101101110001011011000111101110111110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110101111100100111110111111111010110111111101001111011101101100111111011110010111111111100111100101110101101111111010111111110111010110100011111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111010111011111111111100101100111111111111111100111011111111101110110110111010100010100111111110010110110111111100110010111111011111111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111001110111111111110001111011100010110011101111110101100111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101111101110101111001111000100011110100100100101100110111011111101111011100111111100111111011011011101001011011111101111010011011001111011111111011111111111000100111011111010110011101111011011111111111111000001011110100001111101111111111110010111100011111111110010110101011100110110111101110111000110101101001101111111110111111101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01100011101101110111101011111111001110011111111110011111011101110110010110111111111011100111011111110101100101111111111011110110110111001111110111111011110110010110111001100010110101010110101101011111111011101001100101111101011110011101111011101000010111110111110011010111110111011111111110011011101111111011111111010011101010111100111101100111010101101111000111111011011101111111100111111111111000011001000101001101111110111011100011111101111011111011111001111101111110111011010111111101111111110100001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001110010110011101111110101110111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101110101111101111001111000101011110100100100101100110111011111101111011100111111100111111011011011101011011011111101111010011011101111011111111011111101111000100111011111010110011101111011011111111111111000001011110110001111101111110111110010111100011111111110010010101011100110110111100110111100110101101001101111111110111011101110111001101100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011100111011111011110110010110101111101111111111110111111010101111001110111110101011001111101111010111111111110101101111111010011101101101111111011000010111010000101011111001111101111000110111101101101110011000011011111111111111001010110111101010011110111011111101111111111001101011011101101011100001111111101111111011110111111101101010101111111011101011111101111111101111111111111111011011111101111111101110111101101110001111011100111101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101001011110100111111110111111111011001100101111111111000111011001111101111010111011110001101111110110111110111110001100101111111000111111000111100111111111111110111111111011111111101101111101100111111101111011101110010111111111110111111111110101110111101111111011111010111111111111100101111111101111001001010111101111111011010111111111111110110001100110011001111011111111111101000111101111110000100111111100110011111011101111111111110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111011110010110011101111110101110111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101110101111101111001111000101011110100100100101100110111011111101111011100111111100111111011011011101011011011111101111010011011101111011111111010111101111000100111011111010110011101111011011111111111111000001011110110001111101111110111110010111100011111111110010010101011100110110111100110111100110101101001101111111110111011101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01100011101101110111101011111111001110011111111110011111010101110110010010111111111011100111111111110101100101111111111011110110110111001111111111111011110110110110111001100010110101010110101101011111111011101001100101111101011110011101111011101000010111110111110011010111110111011111111110011011101011111011111111010011101010111100111101100111010101101111000111111011011101111111110111111111111010011001100101001101111110111011100011111111111011101011111011111101111110111011010111111101111111110110001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110110011111011110110010110101111111111111111111111111010101111111111111110101011001111101111010111111111110101101111111110011101101111111111011000010111010000101011111011111111111010110111101101111110010110011011111111111111001011110111101110111100011011111101111111111001101011011111101011100001111111101011111011110111111101101010101111111011111011111101111110101111111111111111010001111101111111001110111101101110001111011100111101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10110110111010110110111011011111110011101110111111110010111111011010100010011111111110111100101001011101010111111111101111111111011111110011010001010011111110011101011111101100011101000111111110111011111110111010111110101101101100100111111011111111110101111111011001111101111111111011001111011111111111111010110011111111111101001000100011100101101001001011101111001110110100111111111011111110011000111100100111111111011000111110000011110111111111011011001001110111111110111011011110011111110101111111010110001111";cor_in <= "11011100011101001011111010100001001101000101001010111010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "01100001101101110111101011111111001110111111111110011111010101111110010110111111111011100111010111110101100101111111111011110110110111001111110111111011110110110110111001100010110101010110101101011111111011101001100101111101011110011101111011101000010111110111110011010111110111011111111110011011101111111011111011010011101010111100111101100111010101101111000111111011011101111111100111111111111000011001100101001101111110111011100011111101111011101011111011111100111110111011010111111101111111110100001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11101001101101110111111111101111001110011111111110011111011101111110110010111111111111100111111111110100101101111111111011110011110111001111101111111011110110110110111001110010110101110110011101111111111001101001100101111101011110011001111111110100110111100111110011010111110110011111111110011011101011111011011011010011101110111100111101100111011111101111010111111011111111111111110111111111111010011001100111001101111111111011100011111111111011101011111111111100111111111011011111111101111111110111000111101101";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111110111011001101101011110111000111010011111100111010101011110001111111110110111110111110101100111111111100111111000111100111111101111110111110111011111111101101111101100111111101111011101110010111111111100111111111110101111111101111111011111010111111111011000101111111011111001001010111001111111011110111110111110110110001100110011001111011111110111101000111101111110000100111111100111011011011101111101010110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010111010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111010101111100111111110111111111010110111111001001111011111101100111011011110010111111111100111110101110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111111100111011111111101110110110111010100010100111111110010110110111111100110010111011011111111001010011110101110011101110111111001010100110011010111111111011111001101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11110111110111111001110111111011001110111111111111111111111111111111011110001111011011101011001011111100111011011111111100101111111101111010001111011101011111100011111101111010111111101000111111011101010101111111101001011010111011111101111001111001001101111010110111111100111011101101111011101111101111011111111011111110110011111110001101011111001111111111101111011101111111110111011011111111111101111111011110100110110111100010111111111111011111111010111111110011111111011111111011111011111101111111001101101110";cor_in <= "11000000100010111011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110011010110111011111011110110011110111111101111111111110111111010101111001110111110101011001111101111010111111111110101101111111010011101101101111111011000010111010000101011111001111101111000110111101101101111011110011011111111111111001010110111101110111101111010111101111111111001101011011101101011110001011111101011111011110111111001101010101111111011111011111101111111101111111111111111011001111101111110001110111101101110001111011000011101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111111111111001110111111111110011111011101111110010110111111111011100111011111110101101101111111111011110110110111001011101111111011110110110110111001100010110101010110101101011111111011101001100101111101111110011101111011101000010111100111110011010111110111011111111110011011101111111011111011010011101110111100111101100111010111101111000111111011011111111111110111111111111000011001100101001111111110111011100011111111011011101011111011111101111111111011010111111101111111111111001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11101111011110011111011110011111111101101011110100111111111111111111011001101101011111111000111011001111101111010110011110001101111110110111110111110001100111111111100111111000111100111111111111110111111111011111111101101111101100111111111111011101111010111111111110111111111111101110111111111111011111010111111111011100101111111111111001001010111111111111011010011111111111110110001100110011011111011111111110101000111101111110000100111111100111011111011101111101010110111010111101100111010111111111111001110111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10100110100111111011111101101010101111100111111110111111111010110111111000001111011111101100111011011111010111111111100011110100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110011010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111101100111011111101101110110110111010100010100111111110010110110111111101110010111011011111111001010011110101110111101110111111001010100110011010111111111011111001101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111101011101010101100101111100100110111111001110100110111111000101110110111111101100110111101111011111101101011101110000010010111101110010101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111000111110101110111101001111111011011100111011001110101110110111111100110111110101011011100111110111111011111000111110110101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101101101111100100110111111001110100110011111000101110110111111101100110111101111111111101101011101111000010010111101110011101110111011110011111011111010111111100101101101011101011110101011011101011111111000111111011111000111110101110111101001111111011011100111011001110101110110101111100110111110111111011110111110111111011111000111110100101111111111111101011111110011010111011111111111101011001111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101011111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101100101111100100110111111101110100110111111000101110110111111101100110111101111111111101101011101111001010010111101110011101110111011110111111011111011111111100101101101011101011110101011011101011111111000111111011100000111110101110111101011111111011011000111011001110101110110101111100110111110111111111110111111111111011111000111110100101111111111111101011111110011110111111111111111101011011111010010011111110111110111111100101111111101010111111100111111111111110111011110110110101111111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11110111110111111001110111111011001110111111111111111111111111111111011110001111011011101011001011101110111011111111111100101111011101111010001111101001011111100011111101111010111111101000111111011101010101111111101001011010111011111101111001111001001111111010110111111100101011101101111011101111101111011111111011111110110011111110001101011111001111111111101111011101111111110111011011111111111101111111011110100110110111100010111111111111011111111011111111110011111111011111111001111011111101111111001101101110";cor_in <= "11000000100010111011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110110011111011110110010110111111111111111111110111111010101111001110111110101011001111101111010111111111110101101111111010011101101101111111011000010111010000101011111011111101111000110111101101101110011110011011111111111111001010110111101110011100111010111101111111111001101011011111101011100001011111101011111011110111111101101010101111111011101011111101111111101111111111111111010001111101111111001110111101101110001111011100111101110110110101111111110110101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001110010110011101111110101100111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101111101111101111001111000100011110100100100100100110111011111101111011100111111100111111011011011101000011011111101111010011011101111011111111010111111111000100111011111010110011101111011011111111111111000001011110110001111101111110111110010111100011111111110010010101011100110110111100110111000110101101001101111111110111011101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111110111011001101101011110111000111010011111100111010101011110001111111110110111110111110101100111111111100111111000111100111111101111110111111111011111111101101111101100111111101111011101110010111111111110111111111110101110111101111111011111010111111111011000101111111111111001001010111001111111011010111111111111110110001100110011001111011111111111101000111101111110000100111111100111011011011101111101010110111010111111100111010111111101111011110111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101100101111100100110111111001110100110111111000101110110111111101100110111101111011111101101011101110000010010111101110011101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111000111110101110111111001111111011011000111011001110101110110111111100110111110101111011100111110111111011111000111110100101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001110011110011101111110001110111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101110101111101111001111000101011110100100100101100110110011111101111011100111111100111111011011011101010011011111101111010011011101111011111111010111101111000100111011111010100011101111011011111111111111000001011110110001111101111110111110010111100011111111110010010101011100110110111100110111100110101101001101111111110111011101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111111111111001110111111111110011111011101111110010110111111111011100111011111110101101101111111111011110110110111001011101111111011110110110010111001100010110101010110101101011111111011101001100101111101111110011101111011101000010111110111110011010111110111011111111110011011101111111011111011010011101110111100111101100111010111101111100111111011011111111111110111111111111000011001100111001111111110111011100011111101011011101011111011111101111111101011010111111101111111111110001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011110110011111011110110010110111111111111111111110011111010101111011110111110101011001111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111111111010110111101101101110011110011011111111111111001010110111101110111110111010111101101111111001101011011111101011100001111111101011111011110111111101101010101111111011111011111101111111101111111111111111010001111101111110101110111101101010001111011100111101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01101001101101110111111111101111001110011111111110011111011101111110110010111111111111100111111111110100101101111111111011110110110111001111101111111011110110110110111001100010110101010110101101011111111011101001100101111101011110011001111011101000110111100111110011010111110110011111111110011010101011111011111011010011101110111100111101100111010111101111000111111011111111111111110111111111111010011001100111001111111110111011100011111111111011101011111010111100111111111011010111111101111111110110000111101101";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11111111111011110011010110011111111111110001111011101110011111110111111111111001111111111111111101100101111111011110011111100111111111011111111101111110111111111011100111100011011110010101011111110110011111010010010010110100111111100101111111111011110111111000100111110001101101011010110101010111111100011111111111111111110110011110101111100101100111110100101100111101111100111110100011100101011011111010001101110101010111011101110111110110111011111111111010101111101111010101101111011000100010010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111001101010101100101111100100110111111001110100110111111000101110110111111101100110111101111111111101101011101110000010010111101110011101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111000111110101110111101001111111011011000111011001110101110110111111100110111110111111011100111110111111011111000111110100101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101011111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01111111111011110011011110011111111111110001111011101010011110110111111111111001111111111111101101100101111111011110011111100111111111011111111101111110111111111011100111100011011110010101011111110110011111010010010010110100111111100101111111111011110111111000100111110001101101011010110101010111111000011111111111111111111110011110101111100101100111110100101100111100111100111110100011100001011011111010001101110101010111011101110111110110111011111111111010101111101111010101001111011000100010010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111111111011011110111101111111110111111011101000011110111111111111111111111111011111111101110111111110111111101111100111111111111101111111011110111111111111111111110111111110111101011111110111011111111110010011110101111111101101111111111111111011111100100111111011111111011001110101010011111100011111010111111111111111111111101111111111110111110110111111111101111111111111100111110101111111111110111101111101000111011101111111110110111111111111111110111111101111110101101111011000110110011110111111111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110111011111011110110010110111111111111110111111011111010101111011111111110101011101111101111010111111111110101101111111110011111111101111111011000010111010000101011111001111111111010110111101101111110010010011011111111111110001011110111101010111110111010111101101111111001100011011111101011110001111111101111111011110111111001101011101111111011111011111101111111101111111111111111010001111101111110001110111101101110001111011000111101110111110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101101101111100100111111111101110100110011111000101110110111111101110110111101111111011100101011101111000010010111101110011101110111011110011111011111011111111100101101111011101011100101111011111011111111000111111011111000111110101110111101011111111011010100111011001110101110110101111100110111110111111111110111111111111011111000111110100101111111111111101011111110011110111111111111111101011011111010010011111110111110111111100101110111111110111111100111111111111110111011110110110101011111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110111011111011111110010110111111111111111111111011111010101111011111111110101011101111101111010111111111110101101111111110011101111101111111011000010111010000101011111001111111111010110111101101111110011110011111111111111110001010110111101110111110111010111101101111111001101011011111101011110001111111101111111011110111111001101011101111111011111011111101111111101111111111111111000001111101111110001110111101101110001111011000111101110111110101111111110110101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01111111111011110011011110011111111111110001111011101010011110110111111111111001111110111111101101100101111111011110011111100111111111011111111111111111111111111001100111100011011110010101111111110111011111010010011010110100111111100101101111111011110111111000100111110001101111011011110101010111111101011111111111111011011110011110100111100101110101110100101100111100111100111110100011100001011011111010001101110101010111011101110111111110111011011111111010111111101111010101011111011000100110010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111101011101010101100101111100100010111111001110100110111111000101110110111111101100111111101111011111100101111101110000010010111101110010101110111011110011111011111010111111100101101101011101011110101011011101011101111000111111011111000111111101110111111001111111011011100111011001110101110110111111100110111110101011011100111111111111011111000111110110101111111111111101011111110011010111011111111111101011001111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101001101101110111111111101111001110111111111110011111011101111110110110111111111011100111111111110100101101111111111011110110110111001111101111111011110110110110111001100010110101010110111101011111111011101001100101111101011110011001111011101000110111100111110011010111110111011111111110011010101111111011111011010011101110111100111101100111010111101111000111111011111111111111110111111111111010011001100111001111111110111011100011111111011011101011111010111100111111111011010111111101111111110111001111101101";cor_in <= "11000000011101001011111010100001001101000101001011101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "01111111111011110011010110011111111111110001111011101010011111110111111111111001111110111111101101110101111111011110011111100111111111011111111101111110111111111011100111100011011110010101011111110111011011010010010010110100111111100101101111111011110111111000100111110001101111011010110101010111111100011111111111111111010110011110100111100101100101110100101100111100111100111110100011100001011011111010001101110101010111011101110111110110111011011111111010111111101111010101011111011000100010010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11100110100111111011111101111010101111100111111110111111111010110111111001001111011111101100111011011110010111111111100111110100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111111101111111110111111101101111011111100110111011111000111011111111111100101100111111110111101100111011111101101110110110111010100010100111111110010110110111111100110010111011011111111001010011110101110111101110111111001010100110011010111111111011111001101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111110111011111011111011010111110011101110111111110011111111011010100011011111111111111100101010011111011111111111101110111111001011110001010001010011111110011111011111111100011111000111111110111011111111110011111101111101101100110111111011111111110111111111011001111101111111111111101111011111111110111010110011111111111101001010100011100101101011101011101111001111111100111111111011111111011000111110100111111111011010101110100111110111011111111011001011110111111110111011111110011111111101111111010110001111";cor_in <= "11000000011101001011111010100001001101000101001010111010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111010101111111011111111111011101111111111111101111111111110110110110111101111110101111011101110011011101110101111111110111001110111001111101011110011011111111010011111111111110110011000111111111110111111111110111111111111111111101101111111000111111111110111111011111101110110111111011110111111111111111110101010111011111111101111011111011110111111001111110111101011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111111111111111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000101110001000111110" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101101011110100111111110111111111011001100101011111111000111011001111101111010110011110001101111110110111110111110001100101111111100111111000111100111111111111110111110111011111111101101111101100111111101111011101111010111111111110111111111111101110111111111101011111010111111111111100101111111111111001001011111111111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100111011111011101111111010110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110101111100101111110111111111010110111111001001111011101101100111111011110010111111111100111100101110101101111111010111111110111010110100111111101110000111111010111101111101010110111110001010111000111000101111011110111011001111111101111111110111111101101111011111100110111011111010111011110111111100101110111111111111111100111011111111101110110110111010100010100111111110010110110111111100110010111011011011111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011110111011111011111110010110111111111111111111111111111010101111011111111110101011101111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111111111010110111101101101110011110011011111111111111001010110111101110111110111010111101101111111001101011011111101011110001111111101111111011110111111001101010101111111011111011111101111111101111111111111111010001111101111110001110111101101110001111011000111101110110110101111111110110101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111101011101010101101101111100100110111111001110100110111111000101110110111111101110110111101111011111101101011101111000010010111101110011101110111011110011111011111011111111100101101111011101011110101011011101011101111000111111011111100111110101110111101001111111011011100111011001110101110110111111100110111110111111011100111110111111011111000111110100101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101011111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01111111111011110011011110011111111111110001111011101010011111110111111111111001111111111111111101100101111111011110011111100111111111011111111101111110111111111011100111100011011110010101011111110111011111010010010010110100111111100101101111111111111111111000100111110001101111011000110101010111111101011111111111111111011110011110101111100101100111110100101100111100111100111110100011100001011011111010001101110101010111011101110111110110111011111111111010101111101111010101011111011000100010010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111010101111100111111111111111111010110111111001001111011111101100111011011110010111111111100111100101110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111111100111011111101101110110110111010100010100111111110010110110111111100110010111011011111111001010011110101110011101110111111001010100110011010111111111011111001101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111101001101010101100101111100100110111111001110100110111111000101110110111111101100111111101111011111101101011101110000010010111101110010101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111000111110101110111101001111111011011100111011001110101110110111111100110111110101011011100111110111110011111000111110100101111111111111101011111110011010111011111111111101011001111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011101111111110011011110111111111111111011011011101001111110111111111111111001111111011111111101100111111111110111001111100111111111111111111111111110111111111111100111100111001111010101011111110110011111111010010111110100111111100101111111111111111011111000110111110011111101011000110101010011111000011111111111111111111111011110101111101101100111110100101101111101111101111111100111100101011111111110001101110111010111011101110111110110111011111111111010101111101111010101101111011011110010011110111011111110";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011110111011111011110110010110111111111111111111111111111010101111001110111110101011001111101111010111111111110101101111111010011101101101111111011000010111010000101011111001111111111000110111101101101111011110011011111111111111001010110111101110111110111010111101111111111001101011011101101011100001111111101011111011110111111101101010101111111011111011111101111111101111111111111111010001111101111111001110111101101110001111011000111101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11100001101101110111111111101111001110111111111110011111011101111110110110111111111011100111111111110101101101111111111011110110110111001111101111011011110110110110111001100010110101010110111101011111111011101001100101111101010110011001111011101000010111100111110011010111110111011111111110011011101011111011111011010011101110111100111101100111010111101111000111111011111111111111110111111111111010011001100101001111111110111011100011111111011011101011111010111100111111111011010111111101111111110111001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111011101111111011111111111011100111111111111101111111111110110110110111101111110101111011101111011011101110101111111110111001110111001111101011110011011111111010011111111111110110011000111111111111111111111110111111111111111111101101111111000111111111111111111011111101110110111111001110111111111111111110111010111011111111101111011111011110111111001111110111101011011111111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111111110111111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000101110001000111110" ; wait for 10 ns; 
inp_feat <= "10101011011110011111011110011111111101101011110100111111110111111111011001101101011111111000111011001111101111010100011110001101111110110111110111110001100111111111100111111000111100111111101111110111110111011111111101101111101100111111101111011101111010111111111110111111111110101110111101111111011111010111111111111100101111111111111001001010111001111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100111011111011101111101011110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10101111111110011111011110011111111101001111110100111111111111111111011011100101011111111000111111001111101111010110011110001101111110110111110111110001000101111111000111111000111100111111111111110111111111011111111101101111101110111111001110011111111010111111111110111111110110101110111111111101011111010111111111111100101111111101111001001010111111111111011000111111111111110110011100110011011111011111111111101000111101111110100100111101100111011111011111111111011110111010111101100111010111111101111101110111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001100010110001111111110101100111111100011111101111010111010011110001111100010111101110011101001101100111111001111100111111111101111101111101111001111000100011110100000110101100110111011111101111011100111111110111111011011011101011011011111101111010011111101111011110111010111111111010100111011111011110011101111011011111111111111000001011110110001111101111110111110010111000011111111110010010101011100111110111110110111000110101101001101111111110111011101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111110111011111011010111110011101010111111110011111111011010100011011111111111111110101011011111011111111111101110111101001011110011010001010011111110011111011111101100011111011111111110111011111111111011111101111001101100110111111011111111110111111111011001111101111111111110101111111111111110111010111011111111111101001010100011100101101010101011101011101111100100111111111011111111011100111110100111111111111010101110000111110111011111111011001011010111111111111011111110011111111101111111010110001111";cor_in <= "11011000011101001011111010100001001101000101001010111010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111111111011111011010111110011101110111111110011111101011010100011011111111111111110101011011111011111111111101110111101011011110011010001010011111110011111011111111100011111011111111110101011111111111011111101111001101100110111111011111111110111111111011011111101111111111110101111011111111110111010111011111111111101001010100011100101101010101011101111111111100100111111111011111110011100111110101111111111111010101110000111110111011111111011001011100111111111111011111110011111111101111111010111001111";cor_in <= "11000000011101001011111010100001001101000101001010101010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111011110010110011101111110001100111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101111101111101111001111000100011110100100100100100110111011111101111011100111111100111111011011011101000011011111101111010011011101111011111111010111111111000100111011111010110011101111011011111111111111000001011110100001111101111110111110010111100011111111110010010101011100110110111100110111000110101101001101111111110111011101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101101110101111100101111110111111111010110111111001001111011101101100111111011110010111111111100111100101110111101111111010111111110111010110100111111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111010111011111111111100101100111111111111111100111011111111101110110110111010100010100111111110010110110111111000110010111111011111111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111111111011001101101011111111000111010011111100111010101011110001101111110110111110111110101100111111111100111111000111100111111111111110111111111011111111101101111101100111111101111011101110010111111111100111111111111101110111111111111011111010111111111011000101111111101111001001010111101111011011010111110111111110110001100110011001111011111110111101000111101111110000100111101100110011011011101111101010110111010111101100111010111111101111011100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111110111011001101101011110111000111010011111100111010101011110001111111110110111110111110101100111111111000111111000111100111111101111110111110111011111111101101111101100111111101111011101110010111111111100111111111110101111111111111111011111010111111111011000101111111111111001001010111001111111011110111110111111110110001100110011001111011111110111101000111101111110000100111111100111011011011101111101010110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111011111011111011010111110011101110111111110011111111011010100011011111111111111100101010011111011111111111101110111111001011110011010001010011111110011111011111111100011111000111111110111011111111111011111101111101101100110111111011111111110111111111011001111101111111111111101111011111111111111010110011111111111101001010100011100101101011001011101111101110110100111111111011111110011000111110100111111111011010101110100111110111011111111011001011110111111110111011111110011111111101111111010111001111";cor_in <= "11000000011101001011111010100001001101000101001010111010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "11101001101101110111111111101111001110111111111110011111011101111110110110111111111011100111111111110101101101111111111111110110110111001111101111011011110110110110111001100010110111010110111101011111111011101001100101111101010110011001111011101000010111100111110011010111110111011111111110011011101111111011111011010011101111111100111101100111010111101111000111111011111111111111110111111111111000011001110111101111111110111011100011111111011011111011111010111101111111111011010111111101111111110111001111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "00111111101001101010101100101111100100110111111001110100110111111000101110110111111101100110111101111111111101101011101110000010010111101110010101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011101000111110101110111101001111111011011000111011001110101110110111111100110111110101011011100111110111111011111000111110100101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101011111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111001001011110100111111110111111111011001101101011111111000111010011111101111010111011110001101111110110111110111110001100111111111000111111000111100111111111111110111111111011111111101101111101100111111101111011101110010111111111110111111111110101110111111111111011111010111111111011000101111111111111001001010111001111111011010111111111111110110001100110011001111011111111111101000111101111110000100111111100111011011011101111101010110111010111111100111010111111101111011100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011100100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111101101100111100111011111110110010101111111011111111111011100011111111111100111111111110110110110111101111110101111011100111011011101110101111111110111001110111101111101011110011011111111010011110111111110110001000111111101110111111101110111111111111111111101101111111000111111111110111111011111101110110111111001110111111111111111110111010111011111111101111011111011110111111001111110111101011011110101011000111101111011101101110111011111110101101111101111011111101111111111111101111111111011110111111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000101110001000111110" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101111110100111111110111110111011001101101011110111000111010011111100111010101011110001111111111110111110111110001100111111111000111111000111100111111101111110111110111011111111101101111101100111111101111011101110010111111111100111111111110101110111101111111011111010111111111011000101111111001111001001010111001111111011110111111111111110110001100110011001111011111110111101000111101111110000100111101100111011011011101111101011110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111011111011111011010111110011101110111111110011111111011010100011011111111111111100101011011111011111111111101110111111001011110011010001010011111110011111011111111100011111000111111110111011111111110011111101111101101100110111111011111111110111111111011001111101111111111111101111011111111110111010110011111111111101001010100011100101101011001011101111101111110100111111111011111111011000111110100111111111011010101110100111110111011111111011001011110111111110111011111110011111111101111111010110001111";cor_in <= "11000000011101001011111010100001001101000101001010111010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101101110101111100101111110111111111010110111111001001111011111101100111111011110010111111111100111100101110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111111111111100111011111111101110110110111010100010101111111110010110110111111000110010111011011111111001010011110101110011101110111111001010100110011010111111111011111101101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111010011011100001111101111001010000111111111011110110010110101111100111111111110111111010101111101110111010101011001111111111110111011111110100101111111010011101101101111111101000010111010000101011110011111101111001110111101101101110011010011011111111111011001010111111101010011110111011111101111111111001101011011101101011100001011111101011101011111111111101111010100111111011101001111101110111101111111111111111011011111101011101101110111001101010001111011100011101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101101101111100100110111111001110100110011111000101110110111111101110110111101111011111101101011101111000010010111101110011101110111011110011111011111011111111100101101111011101011110101011011111011111111000111111011111100111110101110111101001111111011011100111011001110101110110101111100110111110111111011110111111111111011111000111110100101111111111111101011111110011110111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101011111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111111111011001101101011111111000111010011111101111010101011110001101111110110111110111110001100111111111100111111000111100111111101111110111110111011111111101101111101100111111101111011101110010111111111100111111111110101110111101111111011111010111111111011000101111111111111001001010111001111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100111011011011101111101010110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001110010110011101111110101100111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101110101111101111001111000101011110100100100101100110111011111101111011100111111100111111011011011101010011011111101111010011011101111011111111011111101111000100111011111010110011111101011011111111111111000001011110110001111101111110111110010111100011111111110010010101011100110110111100110111100110101101001101111111110111011101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01111111111011110011010110011111111111110001111011101010011110110111111111111001111110111111101101110101111111011110011111100111111111011111111111111110111111111001100111100011011111010101011111110110011111010010010010110100111111100101111111111011111111111000100111110001101111011011110101010111111001011111111111111111011110011110101111100101110101110100101100111100111100111110100011100101011011111010001101110101010111011101110111110110111011011111111010101111101111010101011111011000100110010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10101011011110011111011110011111111101001111110100111111110111111111011001101101011111111000111011011111101111010101011110001101111110110111110111110001100101111111100111111000111100111111111111110111111111011111111101101111101100111111101111011101111010111111111110111111111110101110111101111111011111010111111111011000101111111101111001001010111101111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100111011111011101111101010110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101111011110011111011110011111111111101111110100111111110111111111011001100101011111111000111011011111101111010100011110001101111110111111110111111001100101111111100111111000111100111111111111110111111111011111111101101111111100111111101111011101111010111111111100111111111111101110111101111101011111010111111111011000101111111101111001001011111111111111011010111111111111110110001100110011001111011111111111101100111101111110000100111101100110011111011101111111011110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111011110010110011101111110101100111101100011111101111010111010011110001101100010111101110011101001101100111111001111100111111111101111101111101111001111000101011110100100100100100110111011111101111011100111111100111111011011011101011011011111101111010011011101111011111111011111111111000100111011111010110011111101011011111111111111000001011110100001111101111110111110010111100011111111110010010101011100110110111101110111100110101101001101111111110111111101110111001100100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111111111011111011110110111001101010011111110011111101001011100011011111111111111111101011011111011111111111101110111101001011110011010011010111111110111111111111101100011111011111111110101011101111110011111101111011111101110111111011111111110111111111111011111101011111111110101111011111111110111110111010111111111101001111100011100101101110101011101011111111101100111111111011111111011100110110101111111111111010101110100111110011011111111111001011000111111111011011111111011111111101111111010111101111";cor_in <= "11001000011101001011111010100001001101000101011010101010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "11110111110111111001110111111011001110111111111111111111111111111111011110101111011011101011001011101110111011111111111100101111011101111010001111101101011111100011111101111010111111101000111111011101010101111111101001011010111011111101111001111001001111111010110111111100111011101101111011101111101111011111111011111110110011111110001101011111001111111111101111011101111111110111011011111111111101111111011110100110110111101010111111111111011111111011111111110011111111011111111011111011111101111111001101101110";cor_in <= "11000000100010111011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "00111111111001101010101100101111100100110111111001110100110111111000101110110111111101100111111101111011111100101011101110001010010111101110010101110111011110011111011111011111111100101101101011101011110101011011111011101111000111111011111100111111101110111111001111111011111000111011001110101110110111111100110111110101011011100111110111110011111000111110110101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "11000000011101000100000110100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101101110101111100100111111111101111010110111111101001111011101101100111111011110011111111111101111100101110101101111111010111111111111010110100111111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111010111011111111111110101100111111111111111100111011111111101110110110111110100110100111111110010110110111111101110010111111011110111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11100110100111111011111101101010101111100111111110111111111010110111111001001111011111101100111011011110010111111111100111110100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111101100111011111101101110110110111010100010100111111110010110110111111101110010111011011111111001010011110101110011101110111111001010100110011010111111111011111001101";cor_in <= "11000000011101001011111010100001001101000101001001010101011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11011011111111101110110111111110001111001100010110001101111110001111111111100011111101111010111010011110001111100010111101110011101001101100111111001111100111111111101110101111101111001111000101011110100100100101100110110011111101111011100111111100111111001011111101011011011111101111010011011101111011111111010111101111010100111111111011110011101111011011111111111111100001011110110001111101111111111110010111100011111111110010110101011100111110111110110111100110101101001111111111110111011101110111001101100110";cor_in <= "11000000011101001011111010100001110010110101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111011110011010110011111111111110001011011101010011111110111111111111001111111111111101101100101111111011110011111100111111111011111111101111110111111111011100111100011011110010101011111110110011011010010010010110100111111100101101111111111111111111000100110110001101111011000110101010111111000011111111111111111111110011110101111100101100111110100101100111101111100111110100011100101011011111010001101110101010111011101110111110110111011111111111010101111101111010101101111011000100010010110111011111111";cor_in <= "11000000011101001011111001011110001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "01100001101101110111101111101111001110011111111110011111011101110110110010111111111011100111111111110100100101111111111011110111110111001111101111111011110110110110111001100010110101010110101101111111111011101001100101111101011110011001111011101000010111110111010011010111110110011111111110011011101011111011111011010011101010111100111101100111010101101111010111111011011101111111100111111111111010011001000111001101111111111011100011111101111011101011111011111100111111111011010111111101111111110110000111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011110111011111011111110010110111111111111111111111011111010101111011111111110101011101111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111111111010110111101101101111011110011011111111111110001010110111101010111110111010111101101111111001101011011111101011110001111111101111111011110111111101101010101111111011111011111101111111101111111111111111010001111101111110001110111101101110001111011100111101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110011011110110011111011111110010110111111111111111111111111111010101111011101111110101011101111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111101111010110111101101101110011110011111111111111111001010110111101110111100111010111101111111111001101011011111101011110001011111101011111011110111111001101010101111111011111011111101111111101111111111111111010001111101111110001110111101101010001111011000111101110110110101111111110111101100011111001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111011111011111011010111110011101010111111110011111111011010100011011111111111111110101011011111011111111111101110111101011011110001010001010011111110011111011111111100011111010111111110111011111111110011111101111101101100110111111011111111110111111111011011111101111111111110101111111111111110111010110011111111111101001010100011100101101010101011101111101111111100111111111011111111011000111110101111111111011010101110000111110111011111111011001011110111111110111011111110011111111101111111010111001111";cor_in <= "11000000011101001011111010100001001101000101001010111010100111010001110100111110" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111111101111001110011111111110011111011101111110110010111111111111100111111111110100100101111111111011110111110111001111101111111011110110110110111001100010110101010110101101011111111011101001100101111101011110011001111011101000110111100111110011010111110111011111111110011011101011111011111011010011101110111100111101100111010111101111010111111011011111111111110111111111111010011001100111001111111111111011100011111111011011101011111011111100111111111011010111111101111111110110000111101111";cor_in <= "11000000011101001011111010100001001101000101001010101010011000100001110111000001" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110011011100111011111011110110010100101111111111110011111111111011101111111111111110101011101111101111010111111111110101101111111110111111111111111111011000011111010000101011111001111111111010110111101101111110110110011111111111111111001000110111101110111111011010111101111111111001000011011111101011110001111011101111111011110111111001111011111111111011111011111101111111101011111111111111000101111101111110101110111101101110001011011000111101110111110101111111110111101100011110001";cor_in <= "11000000011101001011111010100001001101001010110110101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11110111110111111001110111111011011110111111111111111111111111111111011111001111011011101011001011101110111011111111111100101111011101111010001111101101011111100011111101111010111111101000111111011101010101111111101001011010111011111101111001111001001101111010110111111100111011101101111011101110111111011111111011111110110011111110001101011111001111111111101111011101111111110111011011111111111101111111011110100110110111100010111111111111011111111010111111110011111111011111111001111011111101111111001101101110";cor_in <= "11000000100010111011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111111101111110100111111110111111111011001100101011111111000111011011111101111010110011110001101111110110111110111110001100111111111100111111000111100111111111111110111111111011111111101101111101100111111101111011101111010111111111110111111110111101110111101111101011111010111111111011000101111111101111001001011111101111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100110011111011101111111010110111010111101100111010111111101111001100111";cor_in <= "00111111011101001011111010100001001101000101001010101010011000100001110100111110" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111011111111111111111111111011101111111011111101111011111110111110111111111011110101111001111111011011101110101111111110111001110111111111101011110011111110111010011111111111110110011010111111111111111111111110111111111111111111101101111111100111111011110111111111111101110110111111011110111111111111111110101010111011111111100111111111111110111111011111110111111111011110111111000111101111011101111110111011111110100111111101111011011101111111111111111111111111111110111111";cor_in <= "11000101010101001011111010100001001101000101001010101010011000101110001000111110" ; wait for 10 ns; 

      -- insert stimulus here 

      wait;
   end process;

END;
