--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:52:57 07/25/2019
-- Design Name:   
-- Module Name:   D:/siva/Masters/Thesis/07_ETE_19/part_svhn/cifat_full_tb.vhd
-- Project Name:  part_svhn
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: cifar_full_check
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY cifat_full_tb IS
END cifat_full_tb;
 
ARCHITECTURE behavior OF cifat_full_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT cifar_full_check
    PORT(
         inp_feat : IN  std_logic_vector(511 downto 0);
         cor_in : IN  std_logic_vector(79 downto 0);
         cor_out : OUT  std_logic_vector(79 downto 0);
         out_fin : OUT  std_logic_vector(79 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal inp_feat : std_logic_vector(511 downto 0) := (others => '0');
   signal cor_in : std_logic_vector(79 downto 0) := (others => '0');

 	--Outputs
   signal cor_out : std_logic_vector(79 downto 0);
   signal out_fin : std_logic_vector(79 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: cifar_full_check PORT MAP (
          inp_feat => inp_feat,
          cor_in => cor_in,
          cor_out => cor_out,
          out_fin => out_fin
        );

   -- Clock process definitions
   --<clock>_process :process
   --begin
		--<clock> <= '0';
		--wait for <clock>_period/2;
		--<clock> <= '1';
		--wait for <clock>_period/2;
   --end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      --wait for <clock>_period*10;
inp_feat <= "01111111111011110011010110011111111111110001111011101010011111110111111111111001111110111111101101100101111111011110011111100111111111011111111111111110111111111001100111100011011110010101111111110111011111010010010010110100111111100101101111111011110111111000100111110001101111011001110101010111111101011111111111111111010110011110100111100101100101110100101100111100111100111110100011100001011011111010001101111101010111011101110111110110111011011111111010111111101111010101011111011000100110010110111011111111";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111111111011110110111011111111110111111111111011101111111111111101111111111110111110111111111011110101111011101111011011101110101111111110111001110111001111101011110011011111111010011111111111110110011010111111111111111111111110111111111111111111101101111011100111111011110111111111111101110110111111011110111111111111111110101010111011111111101111011111011110111111011111110111111011011110111011000111101111011101111110111011111110101111110101111011011101111111111111101111111111111110111111";cor_in <= "10111111101110011100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11111111011101111110111101111011111110111011111111111111111111111011101111111111111101111111111110111110111111111011110101111001111111011011101110101111111110111001110111111111101011110011011111111010011111111111110110011010111111111111111111111110111110111111111111101101111111000111111011110111111111111101110110111111011110111111111111111110101010111011111111101111111111111110111111011111110111111011011110111011000111101111011101111110111011111110100111111101111011011101111111111111111111111111111110111111";cor_in <= "11000001101110011100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11101111011110011111011110011111111101101011110100111111111111111111011001101101111111111001111011001111101111010110011110001101111110110111110111111101101111111111100111111000111100111111111111110111111111011111111101101111101100111111111111011101111010111111111110111111111111101110111111111111011111011111111111011100101111111111111001001010111011111111011010111111111111110110011100110011011111011111111111101100111101111110001100111111100111011111011101111101111110111010111111100111010111111111111011110111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11100110100111111011111101101010101111100111111110111111111010110111111001001111011111101100111011011110010111111111100111100100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111111100111011111101101110110110111010100010100111111110010110110111111100110010111011011111111011010011110101110011101110111111001010100110011010111111111011111001101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110100111100100111111111101111010110111111101001111011101111100111111011110011111111111100111100101110101101110111010111111110111110110100010111101110000111111010111101111101010110111110001010011000111000101111010110111111011111101101111111110111111101101111011111100110111011111010111011111111111110101101111111111111111100111011111011101110110110111110101110101111111110010110110111111001110010111111011110111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111101110111111011110111111101111110111111111111011111111111001111011111001101101001101011011011101110111011111111111100101111011111101000001111001101011111100011111111111010111111101000111111011101111101110111111101011010110111111111111001111101011111111011110111111100111011111101111011101110111111111111111010111111110111111110001101011111001111111111101101011101111111110111011011111110111101111111011110110110111111100010111111111011011111111011111111110011111111011111101001111011111101111111101101100110";cor_in <= "10111111010000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110100111100101111111111101111010110111111101001111011101111100111111011110011111111111101111100101110101100110111010111111111111010110100011111101110000111111010111101111101010111111110001010011000111010101011110110111111001111101101111111110111111101101111011111100110111011111010111011110111111100101110111111111111111100011010111011101110110110111110101110100111111110010110110111011001110010111111011110111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01111111111011110011010110011111111111110001111011101010011111110111111111111001111110111111101101110101111111011110011111100111111111011111111011111110111111111001100111100011011110010101111111110111011111010010010010110100111111100101101111111011110111111000100111110001101111011011110101010111111101011111111111111011011110011110101111100101110101110100101100111100111100111110100011100001011011111010001101110101010111011101110111111110111011011111111010101111101111010101011111011000100110010110111011111111";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11110111110111111001110111111011000110111111111111111111111111111111011111001111101011101011001011101110111011111111111100101111011101111010001111101101011111100011111101111010111111101000111111011101010101111111101101011010111011111101111001111001011111111010110111111100111011101101111011101110101111011111111011111110110011111110001101011111001111111111101101011101111111110111011011111111111101111111011110100110110111100010111111111111011111111011101111110011111111011111111001111011111101111111001101100110";cor_in <= "10111111010000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101001111110100111111110111111111011001101101011111111000111011001111101111010110011110001101111110110111110111110001100101111111100111111000111100111111111111110111111111011111111101101111101100111111101111011101111010111111111110111111111111101110111101111101011111010111111111111100101111111111111001001010111111111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100111011111011101111111011110111010111101100111010111111101111001100111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100011101101110111101011111011001110111111111110011111010101110110010110111110111011100111010111110101100101111111111011110110110111001011110111111011110110010010111101100010110101010110101101010111111011111001100101111101111110011101111011101000010111110111010011010111110111011111111110011011101011111011111111010011101010111100111101100111010101101111100111101011011100111111100111101111111000011001000101001101111110111001100011111101111011101011111001111101111110101011010110111100110111110100001111001111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110110011111011110110010110101111111111111111111111111010101111001111111110101011001111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111101111010110111101101111110010110011011111111111111001010110111101110111100011010111101101111111001101011011111101011100001011111101011111011110111111101111010101111111011111011111101111111101111111111111111010001111101111111001110111101101110001111011100111101110110110101111111110111101100010111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111110111010111011111011011111110011101110111111110011111111011010100010011111111111111100101011011101010111111111101111111111011111110011010001010011111110011101011111111100011101000111111110111011111110111011111100101101101100110111111011111111110101111111011001111101111111111011001111011111111111111010110011111111111101001010100011100101101001001011101111101110110100111111111011111110011000111110100111111111011000101110100011110111111111111011001011110111111110111011111110011111111101111111010110001111";cor_in <= "10111111110000001100000010111010110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111111101111001110111111111110011111011101111110010010111111111011100111111111110101101101111111111011110110110111001111101111111011110110110110111001100010110101010110101101011111111011101001100101111101011110011001111011101000010111100111110011010111110111011111111110011011101111111011111011010011101110111100111101100111010111101111000111111011011111111111100111111111111010011001100101001101111110111011100011111111011011101011111010111100111111111011010111111101111111110110001111101111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11101111011101111111111100111011111110111011111111111111111111111111101011111111111111111111111110110110110111111111110101111001101110011111101110101111111110111101010111111111101011110011011111111010111111111111110110011101111111111110111111101110111110111111111111101101011111000111111111110111111111111101110110111111001110111111111111111010101010111011111111101111111111111110111111011111110111111111011110111111000111101111011101111110111011111110100111111101111011111111111111111111111111111111011110111111";cor_in <= "10110010110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011110110011111011110110010110111111111111111111111111111010101111011100111110101011001111101111010111111111110101101111111110011101101101111111011000010111010000101011111001111101111010110111101101101110011110011111111111111111001010110111101110111110111010111101101111111001101011011111101011110001011111101011111011110111111001101010101111111011111011111101111111101111111111111111000001111101111110001110111101101010001111011000111101110110110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111011111011111011010111110011101110111111110011111111011010100011011111111111111100101011011111011111111111101110111111001011110011010001010011111110011111011111111100011111000111111110111011111111111011111101111101101100110111111011111111110101111111011001111101111111111111101111011111111111111010110011111111111101001010100011100101101011001011101111101111110100111111111011111110011000111110100111111111011010101110100011110111011111111011001011110111111110111011111110011111111101111111010110001111";cor_in <= "10111111110000001100000010111010110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111011111111111011111111111011101111111111111101111111111110110110110111101111110101111011101111011011101110101111111110111001110111001111101011110011011111111010011111111111110110011000111111111111111111111110111111111111111111101101111111000111111111110111111011111101110110111111011110111111111111111110111010111011111111101111011111011110111111001111110111101011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111111110111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11100110100111111011111101111010101111100111111110111111111010110111111001001111011111101100111011011110010111111111110011110101110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111001111000101111011110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111101100111011111101101110110110111010100010100111111110010110110101111101110010111011011011111001010011110101110111101110111111001010100110011010111111111011111001101";cor_in <= "11000000110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111011111011111011010111111011101110011111110011111101011010100011011111111111111111101001011111011111111111101110111111001011110001010011010011111110111111011111100100011111001111111110111011111011111011111101111101101100110111111011111111110111111111011001111101011111111110101111001111111110111010111011111111111101001010100011100101101010101011101011111111100100111111111011111111011100111100101111111111111010101110000111110111011111111011001011010111111111011011111110011111111101111111010110001111";cor_in <= "10110000110000001100000010111010110000001011110110101110010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101001111110100111111110111111111011011101101011111111000111011001111101110010100011110001101111110110111110111110001100101111111000111111000111100111111101111110111110111011111111101101111101100111111101111011101111010111111111110111111111110101110111101111101011111010111111111111100111111111111111001001011111001111111011010111111111111110110011100110011001111011111111111101000111101111110000100111101100111011111011111111111011110111010111101100111010111111101111001100111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011000011111011110111111111110111111001010110110101101111111101111111101100011011101111010111110011110001111100110111101111011101100111100111111001111100111101111101111101110111111111111110100111110100111110111101111111111111101111111100111011100111011011111111101011111011111101111110011111001111111110111111111110111000100111111111011100011111111011011111011111111000111111110101101111111111111111111110110100011111101111110010110011101100111111101110111001110101101111101111011110111011101111111011100100110";cor_in <= "00100000110000001100000010111010001111111011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111011111111001110111111111110011111011101111110010110111111111011100111011111110101100101111111111011110110110111001111101111111011110110110110111001100010110101010110101101011111111011101001100101111101011110011101111011101000010111110111110011010111110111011111111110011011101111111011111111010011101010111100111101100111010101101111000111111011011101111111110111111111111000011001100101001101111110111011100011111111011011101011111011111100111110111011010111111101111111110100001111101111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011100111111111011110110010110101111101111111111110111111010101111001110111110101010001111111111110111111111110100101111111010011101101101111111011000010111010000101011110011111101111000110111101101101111011000011011111111111111001010110111101010011110111011111101111111111001101011011101101011100001111111101011101011110111111101101010101111111011101011111101111111101111111111111111011011111101111111101110111101101110001111011100111101110110110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "00111111101011101010101100101111100100010111111001110100110011111000101110110111111101100111111101111011111100101011101111001010010111101110011101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111100111110101110111101011111111011011100111011001110101110110111111100110111110111111011110111111111111011111000111110100101111111111111101011111110011010111011111111111101011001111010011011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001110010110011101111110001100111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101110101111101111001111000101011110100100100100100110110011111101111011100111111100111111011011011101010011011111101111010011011101111011111111011111111111000100111011111010100011101111011011111111111111000001011110100001111101111110111110010111100011111111110010010101011100110110111100110111000110101101001101111111110111011101110111001100100110";cor_in <= "10111111110000001100000010111010001111111011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "10101011011110011111011110011111111001001011110100111111110111111111011001101101011111111000111011011111101111010101011110001101111110110111110111110001100111111111000111111000111100111111101111110111110111011111111101101111101100111111101111011101111010111111111110111111111110101110111101111111011111010111111111011000101111111111111001001010111001111111011010111111111111110110001100110011001111011111111111101000111101111110000100111101100111011111011101111101011110111010111101100111010111111101111001100111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101001101101110111111111101111001110111111111110011111011101111110110110111111111011100111111111110101101101111111111111111110110111001111101111111011110110110110111001100010110111010110111101011111111011101001100101111101010111011001111011101000010111100111110011010111110111011111111110011010101111111011111011010011101111111110111101100111010111101111000111111011111111111111110111111111111000011001110111101111111110111011101011111111011011111011111010111100111111111011011111111101111111111111001111101100";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101101110101111100101111110111111111010110111111001001111011101101100111111011110010111111111100111100101110111101111111010111111110111010110100111111101110000111111010111101111101010110111110001010111000111000101111010110111011001111111101111111110111111101101111011111100110111011111010111011110111111100101100111111111111111100111011111111101110110110111010100010100111111110010110110111111100110010111011011011111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110100111100100111111111101111010110111111101001111011101101100111011011110011111111111100111100101110101101111111010111111111111110110100011111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111010111011111111111100101100111111111111111100111011111111101110110110111110100110100111111110010110110111111100110010111111011110111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110011011110111011111011110110010110111111111111111111111111111010101111001110111110101011001111101111010111111111110101101111111010011101101101111111011000010111010000101011111001111111111000110111101101101111011110011011111111111111001010110111101110111111111010111101111111111001101011011101101011110001111111101011111011110111111101101010101111111011111011111101111111101111111111111111001011111101111111101110111101101110001111011000111101110110110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011001111111001000111111111111001111011010011111001111111010101101111111110011011101111010111110110111101101100111111101111011101010101100101111001111101111111111101111101110101111011111010100111110101111110101100110111111110101111111110111011111111111011011111101001111011111001101010010011011111011110110011100110111000101111111111010110011101111011011111111111111000111111111100111111101111111111111011110110011101101111011110110010100111111111100111111001110101101001100111011110111111101110111001111111110";cor_in <= "10111111110000001100000010111010001111111111111110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110110011111011110110010110101111111111110011111111111011101111011111111110101011101111101111010111111111110101101111111110011111111101111111011000010111010000101011111001111101111010110111101101111110011010011011111111111110001001110111101110111110011010111101101111111001100011011111101011100001111011101111111011110111111001101011101111111011111011111101111111101111111111111111010101111101111110001110111101101110001111011100111101110111110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100011101101110111101011111111001110011111111110011111010101110110010010111110111011100111010111110101100101111111111011110110110111001111110111111011110110010010111101100010110101010110101101011111111011111001100101111101011110011101111011101000010111110111010011010111110111011111111110011011101011111011111111010011101010111100111101100111010101101111000111111011011100111111100111101111111000011001000101001101111110111011100011111101111011101011111001111101111110111011010111111101111111110100001111101111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101100111111100100110111111101110100110111111010101110111111111101101110111101111111111111101011101111011010010111101110011101110111011110111111011111011111111110101101111011111011110101111011111011111011100111111011101100111110101110111101111111101111011100111011001110101110110101111101110111110111111111110111111111111011111000111110100111111111111111101111111111011111111111111111111101011011110110011011111110111110111101101101111111111011111111100111101111111110111011110110110101111111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011011111111101110110111111110001111001110010110011101111110101111111101100011111101111010111010011110001101100010111101110011101001101100111111001111100111111111101111101111101111001111000101011110100100100101100110110011111101111011100111111100111111011011011101011011011111101111010011011101111011111111011111101111010100111011111011110011101111011011111111111111000001011110110001111101111110111110010111100011111111110010010101011100110110111110110111100110101101001101111111110111011101110111001100100110";cor_in <= "10111111110000001100000010111010001111111011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111110111111001110111111001101110111111111111111111111111001111011111001101101001101011011011101110111011111111111100101111011101111000001111101101011111100011111101111010111111101000111111011101110101110111111101011010111011111111111001111101011111111011110111111100111011111101111011101110111111011111111010111111110111110110001001011111101111111111101101011101111111110111011011111110111101111111011110110110110111100010111111111111011111111011111111110011111111011111101001111011111101111111001111100110";cor_in <= "10111111010000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100011101101110111101111111111001110011111111110011111010101110110010010111110111011100111010111110101100101111111111011110110110111001111110111111011110110010110111001100010110101010110101101011111111011101001100101111101011110011101111011101000010111110111010011010111110111011111111110011011101011111011111111010011101010111100111101100111010101101111010111111011011100111111110111111111111010011001000101001101111111111001100011111101111011101011111001111100111110111011010111111101111111110100001111101111";cor_in <= "10111111110000001100000010111010110000001010110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110011011110111011111011110110011110111111111111111111110111111010101111001110111110101011001111101111010111111111110101101111111010011101101101111111011000010111010000101011111001111101111000110111101101101111011110011011111111111111001010110111101110111111111010111101111111111001101011011101101011110001011111101011111011110111111001101010101111111011111011111101111111101111111111111111011011111101111111101110111101101110001111011001011101110110110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001100010110011101111110101100111101100011111101111010111010011110001101100010111101110011101101101100111111001111100111111111101111101111101111001111000100011110100100110101100110111011111101111011100111111100111111011011011101011011011111101101010011011101111011110111011111101111000100111011111011110011101111011011111111111111000001011110100001111101111111111110010111100011111111110010010101011100111110111100110111000110101101001101111111110111111101110111001100100110";cor_in <= "10111111110000001100000010111010001111111011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110101111100101111111111111111010110111111001001111011101101100111011011110010111111111100111100101110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111011110111011001111101101111111110111111101101111011111100110111011111010111011111111111100101100111111111111111100111011111111101110110110111010100010100111111110010110110111111000110010111111011111111001010011110101110011101110111111001010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110110011111011111110010110111111111111111111111011111011101111011111111110101011101111101111010111111111110101101111111110011111111101111111011000010111010000101011111001111111111010110111101101111110010110011011111111111111001011110111101110111110111010111101101111111001100011011111101011110001111111101111111011110111111001101011101111111011111011111101111111101111111111111111010001111101111110001110111101101110001111011000111101110111110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110101111100111111111111111111010110111111101001111011101101100111011011110010111111111100111100100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111011110111011001111111101111111110111111101101111011111100110111011111000111011111111111100101101111111110111111100111011111111101110110110111010100010100111111110010110110111111100110010111111011111111011010011110101110011101110111111011010100110011011111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111111111011001101101011111111000111010011111100111010101011110001111111110110111110111110001100111111111000111111000111100111111101111110111110111011111111101101111101100111111101111011101110010111111111110111111111110101111111111111111011111010111111111011000101111111111111001001010111001111111011010111111111111110110011100110011001111011111111111101000111101111110000100111111100111011011011101111101010110111010111111100111010111111101111011100111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100011101101110111101011111011001110011111111110011111010101110110010110111110111011100111010111110101100101111111111011110110110111001011110111111011110110010010111101100010110101010110101101010111111011111001100101111101111110011101111011101000010111110111010011010111110111011111111110011011101011111011111111010011101010111100111101100111010101101111100111101011011100111111110111101111111000011001000101001101111110111001100011111101111011101011111001111101111110101011010110111100111111110100001111001111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11111111111111110011010110011111111111110001011011101110011110110111111111111001111111111111111101100111111111011111011111100111111111011111111111111110111111111011100111100011011110010101011111110110011111010010010010110100111111100101111111111111111111111000100111110011101111011000110101010111111100011111111111111111111110011110101111101101100111110100101100111101111101111110100011100101011011111010001101110101010111011101110111110110111011111111111010111111101101010101101111011000110010010110111011111111";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11110100110111111111110111110111011110111111011111111111101111011111011111000101110101101111111011011110111111111010111100111111111111101110101111101000111001101011111101111010111111111010111110011111101111111111111101111111111111011111111011111101011111111011111111111101110011111111111111101111111111111111111101101111111111110111111101111111011111111111111111010111111111111111011111111111111111111111011111101111111111111110111011111111111001111111111111110111111101011111101001111111111101101011111111101110";cor_in <= "10101011010000001100000010111010110000001011110110101110101111101011111100011110" ; wait for 10 ns; 
inp_feat <= "11111110111010111010111011011111110011101110111111110011111111011010100010011111111111111100101011011101010111111111101111111111001111110011010001010011111110011101011111111100011101000111111110111011111110111010111110101101101100100111111011111111110101111111011001111101111111111011001111011111111111111010110011111111111101001010100011100101101001001011101111101110110100111111111011111110011000111110100111111111011000111110000011110111111111111011001011100111111110111011111110011111111101111111010110001111";cor_in <= "10111111110000001100000010111010110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110101111100100111111111111111010110111111101001111011101111100111111011110010111111111110111100101110101101111111010111111110111010110100011111101110000111111010111101111101010110111110001010111000111000101111010110111111001111101101111111110111111101101111011111100110111011111010111011110111111100101110111111111111111100011011111111101110110110111110100110100111111110010110110111011001110010111111011110111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111111101111001110111111111110011111011101111110110010111111111011100111111111110100100101111111111011110110110111001111101111111011110110110110111001100010110101010110101101111111111011101001100101111101011110011001111011101000010111100111110011010111110111011111111110011010101011111011111011010011101110111100111101100111010111101111010111111011011111111111100111111111111010011001100101001101111111111011100011111111011011101011111010111100111111111011010111111101111111110110001111101101";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11111111111101101110111100111011111110111010101111111011111111111011101011111011111101111111111110110110110111101111110101111001100111011011101110101111111110111101010111111111101011110011011111111010011110111111110110011001111111111111111111101110111111111111111111101101111111000111111011110111111011111101110110111111011110111111111111111110101010111011111111101111011111011110111111011111110111111011011110111011000111101111011101100110111011111110100111111101111011011101111111111111111111111111011111111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11011101111111111011011110101111111111111111011011111101111110101111111111111110111111011111111101101011111110111111101111111110111111111111111111111111111111111111111111110111111110011101111011110111011111111111011111110110111011101101111111111111111111101010110111011011111101011010111101010111101001111111111111111111111111111111101111111101110111111100101101111101101111111011111111111101111101111110111101110101110111011111111111110111111111111111111010101111101111110111111111011001111010010110111011111111";cor_in <= "10111111110000001100000000111111110000000010101110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011101111111110011011111111111111111111001011011101101011110111111111111111000100111111111111111110111111111110111101111110111111111111101111111011110111011111111101111100111101111011101011111111110011011110010010110110100111111100101111111111101111111101000110111110011111111011100110101010011111100011111111111111111110110011110101111101011100111110100101111111101111111111111100111110101011111111110011101110101010111011101110111110110111111111111111110101111101101010101101111011001110100011110111111111110";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111011101111111011111111111011101111111111111101111111111110110110110111101111110101111001101111011111101110101111111110111001110111111111101011110011011111111010011111111111110110011000111111111110111111101110111111111111111111101101111111000111111111110111111011111101110110111111011110111111111111111110101010111011111111101111011111011110111111011111110111101011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111011111111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11111111111101101110111101111011111110111010101111110011111111111011100111111111111100111111111110110110110111101111110101111011101111011011101110101111111110111001110111001111101011110011011111111010011110111111110110011000111111111111111111111110111111111111111111101101111111000111111011110111111011111101110110111111011110111111111111111110111010111011111111101111011111011110111111001111110111101011011110111011000111101111011101101110111011111110101111110101111011011101111111111111101111111111111110111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11111111111111111011111011010111110011101110111111110011111101011010100011011111111111111110101011011111011111111111101110111101001011110011010001010011111110011111011111111100011111010111111110101011101111111011111101111001101100110111111011111111110111111111011011111101111111111110101111011111111110111010110011111111111101001010100011100101101111101011101111111111100100111111111011111111011100111110100111111111111010101110100111110011011111111011001011100111111111111011111110011111111101111111010111001111";cor_in <= "10111111110000001100000010111010110000001011110110101100010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111111111011111011010110111011101110011111110011111101001010100011011111111111111111101011111111011111111111101110111101011011110011010011010111111110111111111111101101011111010111111110101011111111111011111101111101101100110111111011111111110111111111111011111101011111111110101111001111111110111110111011111111111101001010100011100101101110101011101011111111100100111111111011111111011100110100101111111111111010101110100111110011011111111011001011000111111111011011111110011111111111111111010111101101";cor_in <= "10111111110000001100000010111011110000001010110110101110010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111111111101011111101110101011111111011111001111111010101111111111111110011111011111011101111011101011110101011101111111111010111111111110101101111101110111101111101111111011000111110010000101011111101111111111010110111101101111110111110011111111111111110001001110111101010111110101010011101101111111001100111111111101011110001111111101111111011110111111111101011111110111011111111111111111111101011111110111111001001111101111110001111111111101111011011011000111101110111101111011111110110011100011111101";cor_in <= "10111111110000001100000010110011110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111100111111011111101101110100111100101111111111101111010111111111101001111011101111111111111011110011111111111101111100101110101101110111010011111111111110111111010111111110010111111010111101111101000110111110001010011000111010101011111110111111011111101101111111110101111101101111011111100110111011111010111011111111111110111101111111111111111100011011111011101110110110111110111110101111111111010110110111111000110010111111011010111011110011110111110111101110111111011010101110011010110111111011111101101";cor_in <= "10111111110000001100000010110011110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "10110110111010111010111011011111110011101110111111110010111111011010100010011111111111111100101011011101010111111111101111111111001111110011010001010011111110011101011111111100011101000111111110111011111110111010111110101101101100100111111011111111110101111111011001111101111111111011001111011111111111111010110011111111111101001010100011100101101001001011101111101110110100111111111011111110011000111110100111111111011000111110010011110111111111111011001011110111111110111011111110011111111101111111010110001111";cor_in <= "10111111110000001100000010111010110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111110111011100001111101110001011110110011111011110110010110111111111111111111111011111010101111011111111110101011101111101111010111111111110101101111111110011101111101111111011000010111010000101011111001111111111010110111101101101110010110011011111111111110001011110111101110111110111010111101101111111001100011011111101011100001111111101111111011110111111101101011101111111011111011111101111111101111111111111111010001111101111110001110111101101110001111011100111101110110110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101111110101111100100111111111111111010110111111101001111011101101100111111011110010111111111100111100101110101101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111010111011111111111100101100111111111111111100111011111111101110110110111110101010100111111110010110110111111001110010111111011110111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111101111111111011111111101111111111111111011111111111101111111111111111101100111111111111011111111111111011011111011111111111111111111111111111111110111011111011111111111111111111111000111111111111011111111011111111110110111011111111111111111101111111111011110111011111111101011001111101010111111101111111111111111111111111111110001111111111111111111100101101111100111111111111101111111111110111111111011101110111110111111111111111111111111111111111111111111111101111011111101111111011111111011010111111111110";cor_in <= "10111111110000001100000000111111110000001010110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101101110101111100101111111111111111010110111111101001111011101101100111111011110010111111111100111100101110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111010111011111111111100101100111111111111111100111011111111101110110110111010100010101111111110010110110111111100110010111011011111111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "00111111101011101010101100101111100100010111111001110100110111111000101110110111111101100110111101111011111100101111101110000010010111101110010101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111100111110101110111101001111111011011100111011001110101110110111111100110111110101011011100111110111111011111000111110110101111111111111101011111110011010111011111111111101011001111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11010111110111111001110111111011001110111111111111111111111111111111011111001111101011101011001011101110111011111111111100101111011101111010001111101101011111101011111101111010111111101000111111011100010101111111111101011010111011111101111001111001011111111011110111111100111011101101111011101110111111011111111010111111110111111110001101011111001111111111101101011101111111110111011011111111111101111111011110100110110111101010111111111111011111111011111111110011111111011111111001111011111101111111001111100110";cor_in <= "10111111010000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101101101111100100110111111001110100110111111000101110110111111101100111111101111011111100101011101110000010010111101110010101110111011110011111011111011111111100101101111011101011110101011011101011111111000111111011111100111110101110111111001111111011011000111011001110101110110111111100110111110101111011100111110111111011111000111110100101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01111111111011110011010110011111111111110001111011101010011111110111111111111001111110111111101101110101111111011110011111100111111111011111111001111110111111111001100111100011011110010101011111110111011011010010010010110100111111100101101111111111111111111001100110110001101111011000110101010111111001011111111111111111010110011110100111100101110101110100101100111100111100111110100011000101011011111010001101111101000111011101110111110110111011011111111010101111101111010101011111011000100110010110111011111111";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111011111011111011010111110011101110111111110011111111011010100011011111111111111100101011011111011111111111101110111111001011110011010001010011111110011111011111111100011111000111111110111011111111111011111101111101101100110111111011111111110111111111011001111101111111111111101111011111111110111010110011111111111101001010100011100101101011001011101111101111110100111111111011111110011000111110100111111111011010101110100111110111011111111011001011110111111110111011111110011111111101111111010110001111";cor_in <= "10111111110000001100000010111010110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111111111101111111101111111111011111111111111110111010101101111111111111011111011111110101111111111011111111111111111111111111111111111110111111111111111111111111111111111111111111111011101111011111111111111111111111111011111110110111111111101111111111111111101111011101111010101111110111111001111110111011110111111111111111011111111111111111111110111111111111111111111011111111111111110111101111111111111111111111111111111110111110111111111101101111101011111111101111111111111110111111110111111111111011";cor_in <= "10111111110000001011011111010100110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11100110100111111011111101101010101111100111111110111111111010110111111001001111011111101100111011011110010111111111100111110100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111101100111011111101101110110110111010100010100111111110010110110111111100110010111011011111111001010011110101110011101110111111001010100110011010111111111011111001101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111010101111111011111111111011100111111111111100111111111110110110110111101111110101111011101111011011101110101111111110111001110111001111101011110011011111111010011111111111110110011000111111111110111111111110111111111111111111101101111111000111111111110111111011111101110110111111011110111111111111111110111010111011111111101111011111011110111111001111110111101011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111011111111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11111111111001101110111101111011111110111010101111110011111111111011100111111111111100111111111110110110110111101111110101111011101111011011101110101111111110111001110111001111101011110011011111111010011110111111110110001000111111101110111111111110111111111111111111101101111111000111111011110111111011111101110110111111011110111111111110111110111010111011111111101111011111011110111111001111110111101011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111011110111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101001011110100111111110111111111011001101101011111111000111011001111101111010110011110001101111110110111110111110101100111111111000111111000111100111111111111110111111111011111111101101111101100111111101111011101111010111111111110111111111111101110111111111111011111010111111111111100101111111111111001001010111001111111011010111111111111110110011100110011001111011111111111101000111101111110000100111111100111011111011101111101111110111010111111100111010111111101111011110111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "00111111101011101010101100101011100100010111111001110100110111111000101110110111111101100111111101111011111101101111101110000010010111111110010101110111011110011111011111011111111100101101101011101011110101011011101011101111000111111011111100111111101110111111001111111011111000111011001110101110110111111100110111110101011011100111110111111011111000111110110111111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "01100001101101110111111111101111001110111111111110011111011101111110110010111111111011100111111111110100100101111111111011110110110111001111111111111011110110110110111001100010110101010110101101111111111011101001100101111101011110011001111011101000010111100111110011010111110111011111111110011011101011111011111011010011101010111100111101100111010111101111000111111011011101111111100111111111111010011001100101001101111111111011100011111111011011101011111010111100111110111011010111111101111111110110001111101111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "11111111111011110011010110011111111111110001111011101010011111110111111111111001111111111111101101100101111111011110011111100111111111011111111111111110111111111011100111100011011111010101111111110110011111010010010010110100111111100101111111111011111111111000100111110001101111011001110101010111111100011111111111111111010110011110101111100101100111110100101100111100111101111110100011100101011011111010001101110101010111011101110111110110111011011111111010111111101111010101001111011000100010010110111011111111";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111011110011011110011111111111110001011011101010011111110111111111111001111111111111101101100111111111011111011111100111111111011111111111111110111111111011100111100011011111010101011111110110011111010010010110110100111111100101111111111011110111111000100111110001101101011010110101010111111000011111111111111111111110011110101111100101100111110100101101111101111100111110100011100101011011111010001101110101010111011101110111110110111011111111111010101111101111010101101111011000100010010110111011111111";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111100111011111110111011101111111011111111111011100011111111111110111111111110110110110111101111110101111011101111011111101110101111111110111001110111111111101011110011011111111010011111111111110110011000111111111110111111101110111111111111111111101101111111000111111111110111111011111101110110111111011110111111111111111110101010111011111111101111111111011110111111001111110111111011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111011111111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111010101111110011111111111011100111111111111100111111111110110110110111101111110101111011101110011011101110101111111110111001110111001111101011110011011111111010011110111111110110011000111111101110111111111110111111111111111111101101111111000111111011111111111011111101110110111111011110111111111111111110111010111011111111101111011111011110111111001111110111101011011110011011000111101111011101101110111011111110101111110001111011011101111111111111111111111111111110111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11110111110111111001110111111001001110111111111111111111111111001111011111001101101011101011001011101110111011111111111100101111011101111000001111101101011111101011111101101010111111101000111111011101110101111111111101011010111011111101111011111101011111111011110111111100111011101101111011101110111111011111111010111111110111111110001001011111101111111111101101011101111111110111011011111110111101111111011110100110110111100010111111111111011111111011111111110011111111011111101001111011111101111111001101100110";cor_in <= "10111111010000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11110111110111110001110111111011001110111111111111011111111111111111011110001111011011101011001011111100111011011111111100101111111111111010001111111001011111100011111101111010111111101000111111011101010111111111101001011010111011011101111001011001001101110010110111111100111011101111111011101111101111011111111011111110110011111110001101011111001111111111101111011001111111011111011011111101111101111101011110100110111011111000111011101111011111111011111111110011111111111111111011111011111101111111001101101110";cor_in <= "10111111010000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111111111011111011010111110011101110111111110011111101011010100011011111111111111111101011011111011111111111101110111101011011110011010011010011111110011111011111111101011111010111111110101011111111111011111101111001101100110111111011111111110111111111011001111101111111111110101111011111111110111010111011111111111101001010100011100101101011101011101111101111100100111111111011111111011100111110101111111111111010101110100111110111011111111011001011010111111111011011111110011111111101111111010111001111";cor_in <= "10111111110000001100000010111010110000001011110110101110010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101101101111100100110111111001110100110011111000101110110111111101110110111101111011111100101011101111000010010111101110011101110111011110011111011111011111111100101101111011101011110101011011101011111111000111111011111100111110101110111101001111111011011100111011001110101110110101111100110111110111111011100111111111111011111000111110110101111111111111101011111110011010111011111111111101011011111010010011111110111110111111100101110111111010111111100111111111111110111011010110110101111111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111110111011100101111101110001011110111011111011111110010100111111111111110111111111111010101111111111111110101011001111101111010111111111110101101111111110011101111101111111011000010111010000101011111001111111111010110111101101101110010110011011111111111110001011110111101010111110111010111101101111111001100011011111101011100001111111101011111011110111111001101011101111111011111011111101111110101011111111111111010001111101111110001110111101101111001111011000111101110111110101111111110111101100011111001";cor_in <= "10111111110000001100000010111010110000000011111010101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "00111111111011101010101101101111100100110111111001110100110011111000101110110111111101110110111101111111111111101011101111001010010111101110011101110111011110111111011111011111111100101101111011101011110101011011101011111111000111111011101100111110101110111101111111111011011100111011001110101110110101111100110111110111111111110111111111111011111000111110100101111111111111101011111110011110111011111111111101011011111010011011111110111110111111100101111111101010111111100111111111111110111011010110110101011111";cor_in <= "10111111110000000100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111010111011111011010111111001101010111111110011111101011010100011011111111111111110101011111111011111111111101110111101001011110001010001010011111111111111011111100100011111011111111110111011111111111011111101111101101100110111111011111111110101111111011011111101111111111110101111011111111110111010110011111111111101001010100011100101101010101011101111111110101100111111111011111110011110111100101111111111111010101110010111110111011111011111001011110111111110011011111110011111110101111111010111001111";cor_in <= "10110011110000001100000011000100110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111001101110111101111011111110111010101111110011111111111011100111111111111100111111111110110110110111101111110111111011101111011011101010101111111110111001110111001111101011110011011111111010011110111111110110001000111111101110111111111110111111111111111111101101111111000111111011111111111011111101110110111111011110101111111110111110111010111011111111101111011111011110111111001111110111101011011110011011000111111111011101101110111011111110101101110001111011011101111111111111111011111111011110111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11100001101101110111111111111111001110111111111110011111011101111110110110111111111011100111011111110101101101111111111011110110110111001111101111011011110110110110111001100010110111010110111101011111111011101001100101111101110111011101111011101000010111100111110011010111110111011111111110011011101111111011111011010011101110111110111101100111010111101111100111111011011111111111110111111111111000011001110101101111111110111011100011111111011011111011111011111100111111111011010111111101111111111111001111101111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111101011111100111111" ; wait for 10 ns; 
inp_feat <= "10100011011110011111011110011111111011101011110100111111110111110111011001101101011110111000111010011111100111010101011110001111111110110111110111110101110111111111000111111000111100111111101111110111110111011111111101101111101100111111101111011101110010111111111100111111111110101111111101111111011111010111111111011000101111111011111001001010111001111111011110111110111110110110001100110011001111011111110111101000111101111110000100111111100111011011011101111101010110111010111111100111010111111101111001100111";cor_in <= "01000000110000001100000010111010110000001011110110110001101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111111110011010110111111111111110001011011101000011110111111111111111001111111111111111101100111111111011111011111100111011101011111111111111110111111111011100111100011011110010101011111111110011111010010010010110100111111100101111111111111111111111000100111110011101111011000110101010111111100011111111111111111110110011110101111101101100111110100101101111101111101111111100111100101011011111010001101110101010111011101110111110110111011111111111010111111101101010101101111011000110010011110111011111110";cor_in <= "10111111110000001100000000111111110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111111111101111110111101111011111110111010101111111011111111111011100111111111111100111111111110110110110111101111110101111011101111011011101110101111111110111001110111001111101011110011011111111010011111111111110110011000111111111110111111111110111111111111111111101101111111000111111111110111111011111101110110111111011110111111111111111110111010111011111111101111011111011110111111001111110111111011011110111011000111101111011101101110111011111110101111111101111011011101111111111111101111111111011110111111";cor_in <= "10111111110000001100000010111010110000001011110110101110101111100110010010111101" ; wait for 10 ns; 
inp_feat <= "11100110100111111011111101101010101111100111111110111111111010110111111001001111011111101100111011011110010111111111100111110100110111101111111010111111110111010110100110111101110000111111010111101111101010110111110001010111000111000101111010110111011001111101101111111110111111101101111011111100110111011111000111011111111111100101100111111110111101100111011111101101110110110111010100010100111111110010110110111111100110010111011011111111011010011110101110011101110111111001010100110011010111111111011111001101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11011011111111101110111111111110001111001110010110011101111110101100111101100011111101111010111010011110001101100010111101110011101001101100111111001111100111111111101111101110101111001111000100011110100100100101100110111011111101111011100111111100111111011011011101011011011111101111010011011101111011111111011111111111000100111011111011110011101111011011111111111111000001011110100001111101111110111110010111100011111111110010010101011100110110111101110111000110101101001101111111110111111101110111001100100110";cor_in <= "10111111110000001100000010111010001111111011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111110100111111011111101100110100111100101111111111101111010101111111101101111011101111100111111011111011111111111101111100101110101101110111010011111011111110111110011111111110000111111011111101111101000111111110001010011000111011111011110110111111001111101101111111110100111101101111011111100110111011111010111011111111111110101111111111111111111100011010111011101110110110111110111110101111111110010110110111011000110010111111011110111011110011110101110111101110111111111010101110011011111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11101110100111111011111101101110101111100101111111111111111010110111111101001111011101101100111111011110010111111111100111100101110111101111111010111111110111010110100111111101110000111111010111101111101010110111110001010111000111000101111011110111011001111111101111111110111111101101111011111100110111011111010111011111111111100101101111111111111111100111011111111101110110110111010100010101111111110010110110111111100110010111111011111111011010011110101110011101110111111011010100110011010111111111011111101101";cor_in <= "10111111110000001100000010111010110000001011110100111100101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101001111110100111111111111111111011001101101011111111000111111001111101111010110011110001101111110110111110111110001100101111111000111111000111100111111111111110111110111011111111101101111101100111111011111011101111010111111111110111111111111101110111111111101011111010111111111111100101111111111111001001010111111111111011000111111111111110110011100110011001111011111111110101000111101111110000100111111100111011111011111111111011110111010111101100111010111111101111101110111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "10101111011110011111011110011111111101101111110100111111110111111111011001101101011111111000111011001111101110010110011110001101111110110111110111110001100111111111100111111000111100111111111111110111110111011111111101101111101100111111101110011101111010111111111110111111110111101110111111111101011111010111111111111100111111111111111001001011111111111111011010111111111111110110011100110011001111011111111111101000111101111110000100111101100111011111011101111111010110111010111101100111010111111101111001100111";cor_in <= "01000000110000001100000010111010110000001011110110101110101111101011111110111101" ; wait for 10 ns; 
inp_feat <= "11111110111010111110111011011111110011101110111111110011111111011010100010011111111111111100101011011101010111111111101111111111001111110011010001010011111110011101011111111100011101000111111110111011111110111010111100101101101100100111111011111111110101111111011001111101111111111011001111011111111111111010110011111111111101001010100011100101101001001011101111101110110100111111111011111110011000111110100111111111011000111110000011110111111111111011001011110111111110111011111110011111110101111111010110001111";cor_in <= "10101111110000001100000010111010110000001011110110110001010000001011111110111101" ; wait for 10 ns; 
      -- insert stimulus here 

      wait;
   end process;

END;
