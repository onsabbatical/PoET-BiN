----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:54:23 07/23/2019 
-- Design Name: 
-- Module Name:    cifar_rinc_40_8 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cifar_rinc_40_8 is
    Port ( inp_feat : in  STD_LOGIC_VECTOR (511 downto 0);
			  cor_out :out STD_LOGIC_VECTOR(79 downto 0);
			  cor_in :in STD_LOGIC_VECTOR(79 downto 0);
           pred_out : out  STD_LOGIC_VECTOR (79 downto 0));
end cifar_rinc_40_8;

architecture Behavioral of cifar_rinc_40_8 is
component LUT8
generic(INIT : std_logic_vector(255 downto 0) := (others => '0') );
port(I0:in std_logic;
I1:in std_logic;
I2:in std_logic;
I3:in std_logic;
I4:in std_logic;
I5:in std_logic;
I6:in std_logic;
I7:in std_logic;
O:out std_logic);
--  Port ( );
end component;
signal C_0_out : std_logic := '0'; 
signal C_1_out : std_logic := '0'; 
signal C_2_out : std_logic := '0'; 
signal C_3_out : std_logic := '0'; 
signal C_4_out : std_logic := '0'; 
signal C_5_out : std_logic := '0'; 
signal C_6_out : std_logic := '0'; 
signal C_7_out : std_logic := '0'; 
signal C_8_out : std_logic := '0'; 
signal C_9_out : std_logic := '0'; 
signal C_10_out : std_logic := '0'; 
signal C_11_out : std_logic := '0'; 
signal C_12_out : std_logic := '0'; 
signal C_13_out : std_logic := '0'; 
signal C_14_out : std_logic := '0'; 
signal C_15_out : std_logic := '0'; 
signal C_16_out : std_logic := '0'; 
signal C_17_out : std_logic := '0'; 
signal C_18_out : std_logic := '0'; 
signal C_19_out : std_logic := '0'; 
signal C_20_out : std_logic := '0'; 
signal C_21_out : std_logic := '0'; 
signal C_22_out : std_logic := '0'; 
signal C_23_out : std_logic := '0'; 
signal C_24_out : std_logic := '0'; 
signal C_25_out : std_logic := '0'; 
signal C_26_out : std_logic := '0'; 
signal C_27_out : std_logic := '0'; 
signal C_28_out : std_logic := '0'; 
signal C_29_out : std_logic := '0'; 
signal C_30_out : std_logic := '0'; 
signal C_31_out : std_logic := '0'; 
signal C_32_out : std_logic := '0'; 
signal C_33_out : std_logic := '0'; 
signal C_34_out : std_logic := '0'; 
signal C_35_out : std_logic := '0'; 
signal C_36_out : std_logic := '0'; 
signal C_37_out : std_logic := '0'; 
signal C_38_out : std_logic := '0'; 
signal C_39_out : std_logic := '0'; 
signal C_40_out : std_logic := '0'; 
signal C_41_out : std_logic := '0'; 
signal C_42_out : std_logic := '0'; 
signal C_43_out : std_logic := '0'; 
signal C_44_out : std_logic := '0'; 
signal C_45_out : std_logic := '0'; 
signal C_46_out : std_logic := '0'; 
signal C_47_out : std_logic := '0'; 
signal C_48_out : std_logic := '0'; 
signal C_49_out : std_logic := '0'; 
signal C_50_out : std_logic := '0'; 
signal C_51_out : std_logic := '0'; 
signal C_52_out : std_logic := '0'; 
signal C_53_out : std_logic := '0'; 
signal C_54_out : std_logic := '0'; 
signal C_55_out : std_logic := '0'; 
signal C_56_out : std_logic := '0'; 
signal C_57_out : std_logic := '0'; 
signal C_58_out : std_logic := '0'; 
signal C_59_out : std_logic := '0'; 
signal C_60_out : std_logic := '0'; 
signal C_61_out : std_logic := '0'; 
signal C_62_out : std_logic := '0'; 
signal C_63_out : std_logic := '0'; 
signal C_64_out : std_logic := '0'; 
signal C_65_out : std_logic := '0'; 
signal C_66_out : std_logic := '0'; 
signal C_67_out : std_logic := '0'; 
signal C_68_out : std_logic := '0'; 
signal C_69_out : std_logic := '0'; 
signal C_70_out : std_logic := '0'; 
signal C_71_out : std_logic := '0'; 
signal C_72_out : std_logic := '0'; 
signal C_73_out : std_logic := '0'; 
signal C_74_out : std_logic := '0'; 
signal C_75_out : std_logic := '0'; 
signal C_76_out : std_logic := '0'; 
signal C_77_out : std_logic := '0'; 
signal C_78_out : std_logic := '0'; 
signal C_79_out : std_logic := '0'; 

signal C_0_S_0_L_0_out : std_logic := '0'; 
signal C_0_S_0_L_1_out : std_logic := '0'; 
signal C_0_S_0_L_2_out : std_logic := '0'; 
signal C_0_S_0_L_3_out : std_logic := '0'; 
signal C_0_S_0_L_4_out : std_logic := '0'; 
signal C_0_S_0_L_5_out : std_logic := '0'; 
signal C_0_S_0_L_6_out : std_logic := '0'; 
signal C_0_S_0_L_7_out : std_logic := '0'; 
signal C_0_S_1_L_0_out : std_logic := '0'; 
signal C_0_S_1_L_1_out : std_logic := '0'; 
signal C_0_S_1_L_2_out : std_logic := '0'; 
signal C_0_S_1_L_3_out : std_logic := '0'; 
signal C_0_S_1_L_4_out : std_logic := '0'; 
signal C_0_S_1_L_5_out : std_logic := '0'; 
signal C_0_S_1_L_6_out : std_logic := '0'; 
signal C_0_S_1_L_7_out : std_logic := '0'; 
signal C_0_S_2_L_0_out : std_logic := '0'; 
signal C_0_S_2_L_1_out : std_logic := '0'; 
signal C_0_S_2_L_2_out : std_logic := '0'; 
signal C_0_S_2_L_3_out : std_logic := '0'; 
signal C_0_S_2_L_4_out : std_logic := '0'; 
signal C_0_S_2_L_5_out : std_logic := '0'; 
signal C_0_S_2_L_6_out : std_logic := '0'; 
signal C_0_S_2_L_7_out : std_logic := '0'; 
signal C_0_S_3_L_0_out : std_logic := '0'; 
signal C_0_S_3_L_1_out : std_logic := '0'; 
signal C_0_S_3_L_2_out : std_logic := '0'; 
signal C_0_S_3_L_3_out : std_logic := '0'; 
signal C_0_S_3_L_4_out : std_logic := '0'; 
signal C_0_S_3_L_5_out : std_logic := '0'; 
signal C_0_S_3_L_6_out : std_logic := '0'; 
signal C_0_S_3_L_7_out : std_logic := '0'; 
signal C_0_S_4_L_0_out : std_logic := '0'; 
signal C_0_S_4_L_1_out : std_logic := '0'; 
signal C_0_S_4_L_2_out : std_logic := '0'; 
signal C_0_S_4_L_3_out : std_logic := '0'; 
signal C_0_S_4_L_4_out : std_logic := '0'; 
signal C_0_S_4_L_5_out : std_logic := '0'; 
signal C_0_S_4_L_6_out : std_logic := '0'; 
signal C_0_S_4_L_7_out : std_logic := '0'; 
signal C_1_S_0_L_0_out : std_logic := '0'; 
signal C_1_S_0_L_1_out : std_logic := '0'; 
signal C_1_S_0_L_2_out : std_logic := '0'; 
signal C_1_S_0_L_3_out : std_logic := '0'; 
signal C_1_S_0_L_4_out : std_logic := '0'; 
signal C_1_S_0_L_5_out : std_logic := '0'; 
signal C_1_S_0_L_6_out : std_logic := '0'; 
signal C_1_S_0_L_7_out : std_logic := '0'; 
signal C_1_S_1_L_0_out : std_logic := '0'; 
signal C_1_S_1_L_1_out : std_logic := '0'; 
signal C_1_S_1_L_2_out : std_logic := '0'; 
signal C_1_S_1_L_3_out : std_logic := '0'; 
signal C_1_S_1_L_4_out : std_logic := '0'; 
signal C_1_S_1_L_5_out : std_logic := '0'; 
signal C_1_S_1_L_6_out : std_logic := '0'; 
signal C_1_S_1_L_7_out : std_logic := '0'; 
signal C_1_S_2_L_0_out : std_logic := '0'; 
signal C_1_S_2_L_1_out : std_logic := '0'; 
signal C_1_S_2_L_2_out : std_logic := '0'; 
signal C_1_S_2_L_3_out : std_logic := '0'; 
signal C_1_S_2_L_4_out : std_logic := '0'; 
signal C_1_S_2_L_5_out : std_logic := '0'; 
signal C_1_S_2_L_6_out : std_logic := '0'; 
signal C_1_S_2_L_7_out : std_logic := '0'; 
signal C_1_S_3_L_0_out : std_logic := '0'; 
signal C_1_S_3_L_1_out : std_logic := '0'; 
signal C_1_S_3_L_2_out : std_logic := '0'; 
signal C_1_S_3_L_3_out : std_logic := '0'; 
signal C_1_S_3_L_4_out : std_logic := '0'; 
signal C_1_S_3_L_5_out : std_logic := '0'; 
signal C_1_S_3_L_6_out : std_logic := '0'; 
signal C_1_S_3_L_7_out : std_logic := '0'; 
signal C_1_S_4_L_0_out : std_logic := '0'; 
signal C_1_S_4_L_1_out : std_logic := '0'; 
signal C_1_S_4_L_2_out : std_logic := '0'; 
signal C_1_S_4_L_3_out : std_logic := '0'; 
signal C_1_S_4_L_4_out : std_logic := '0'; 
signal C_1_S_4_L_5_out : std_logic := '0'; 
signal C_1_S_4_L_6_out : std_logic := '0'; 
signal C_1_S_4_L_7_out : std_logic := '0'; 
signal C_2_S_0_L_0_out : std_logic := '0'; 
signal C_2_S_0_L_1_out : std_logic := '0'; 
signal C_2_S_0_L_2_out : std_logic := '0'; 
signal C_2_S_0_L_3_out : std_logic := '0'; 
signal C_2_S_0_L_4_out : std_logic := '0'; 
signal C_2_S_0_L_5_out : std_logic := '0'; 
signal C_2_S_0_L_6_out : std_logic := '0'; 
signal C_2_S_0_L_7_out : std_logic := '0'; 
signal C_2_S_1_L_0_out : std_logic := '0'; 
signal C_2_S_1_L_1_out : std_logic := '0'; 
signal C_2_S_1_L_2_out : std_logic := '0'; 
signal C_2_S_1_L_3_out : std_logic := '0'; 
signal C_2_S_1_L_4_out : std_logic := '0'; 
signal C_2_S_1_L_5_out : std_logic := '0'; 
signal C_2_S_1_L_6_out : std_logic := '0'; 
signal C_2_S_1_L_7_out : std_logic := '0'; 
signal C_2_S_2_L_0_out : std_logic := '0'; 
signal C_2_S_2_L_1_out : std_logic := '0'; 
signal C_2_S_2_L_2_out : std_logic := '0'; 
signal C_2_S_2_L_3_out : std_logic := '0'; 
signal C_2_S_2_L_4_out : std_logic := '0'; 
signal C_2_S_2_L_5_out : std_logic := '0'; 
signal C_2_S_2_L_6_out : std_logic := '0'; 
signal C_2_S_2_L_7_out : std_logic := '0'; 
signal C_2_S_3_L_0_out : std_logic := '0'; 
signal C_2_S_3_L_1_out : std_logic := '0'; 
signal C_2_S_3_L_2_out : std_logic := '0'; 
signal C_2_S_3_L_3_out : std_logic := '0'; 
signal C_2_S_3_L_4_out : std_logic := '0'; 
signal C_2_S_3_L_5_out : std_logic := '0'; 
signal C_2_S_3_L_6_out : std_logic := '0'; 
signal C_2_S_3_L_7_out : std_logic := '0'; 
signal C_2_S_4_L_0_out : std_logic := '0'; 
signal C_2_S_4_L_1_out : std_logic := '0'; 
signal C_2_S_4_L_2_out : std_logic := '0'; 
signal C_2_S_4_L_3_out : std_logic := '0'; 
signal C_2_S_4_L_4_out : std_logic := '0'; 
signal C_2_S_4_L_5_out : std_logic := '0'; 
signal C_2_S_4_L_6_out : std_logic := '0'; 
signal C_2_S_4_L_7_out : std_logic := '0'; 
signal C_3_S_0_L_0_out : std_logic := '0'; 
signal C_3_S_0_L_1_out : std_logic := '0'; 
signal C_3_S_0_L_2_out : std_logic := '0'; 
signal C_3_S_0_L_3_out : std_logic := '0'; 
signal C_3_S_0_L_4_out : std_logic := '0'; 
signal C_3_S_0_L_5_out : std_logic := '0'; 
signal C_3_S_0_L_6_out : std_logic := '0'; 
signal C_3_S_0_L_7_out : std_logic := '0'; 
signal C_3_S_1_L_0_out : std_logic := '0'; 
signal C_3_S_1_L_1_out : std_logic := '0'; 
signal C_3_S_1_L_2_out : std_logic := '0'; 
signal C_3_S_1_L_3_out : std_logic := '0'; 
signal C_3_S_1_L_4_out : std_logic := '0'; 
signal C_3_S_1_L_5_out : std_logic := '0'; 
signal C_3_S_1_L_6_out : std_logic := '0'; 
signal C_3_S_1_L_7_out : std_logic := '0'; 
signal C_3_S_2_L_0_out : std_logic := '0'; 
signal C_3_S_2_L_1_out : std_logic := '0'; 
signal C_3_S_2_L_2_out : std_logic := '0'; 
signal C_3_S_2_L_3_out : std_logic := '0'; 
signal C_3_S_2_L_4_out : std_logic := '0'; 
signal C_3_S_2_L_5_out : std_logic := '0'; 
signal C_3_S_2_L_6_out : std_logic := '0'; 
signal C_3_S_2_L_7_out : std_logic := '0'; 
signal C_3_S_3_L_0_out : std_logic := '0'; 
signal C_3_S_3_L_1_out : std_logic := '0'; 
signal C_3_S_3_L_2_out : std_logic := '0'; 
signal C_3_S_3_L_3_out : std_logic := '0'; 
signal C_3_S_3_L_4_out : std_logic := '0'; 
signal C_3_S_3_L_5_out : std_logic := '0'; 
signal C_3_S_3_L_6_out : std_logic := '0'; 
signal C_3_S_3_L_7_out : std_logic := '0'; 
signal C_3_S_4_L_0_out : std_logic := '0'; 
signal C_3_S_4_L_1_out : std_logic := '0'; 
signal C_3_S_4_L_2_out : std_logic := '0'; 
signal C_3_S_4_L_3_out : std_logic := '0'; 
signal C_3_S_4_L_4_out : std_logic := '0'; 
signal C_3_S_4_L_5_out : std_logic := '0'; 
signal C_3_S_4_L_6_out : std_logic := '0'; 
signal C_3_S_4_L_7_out : std_logic := '0'; 
signal C_4_S_0_L_0_out : std_logic := '0'; 
signal C_4_S_0_L_1_out : std_logic := '0'; 
signal C_4_S_0_L_2_out : std_logic := '0'; 
signal C_4_S_0_L_3_out : std_logic := '0'; 
signal C_4_S_0_L_4_out : std_logic := '0'; 
signal C_4_S_0_L_5_out : std_logic := '0'; 
signal C_4_S_0_L_6_out : std_logic := '0'; 
signal C_4_S_0_L_7_out : std_logic := '0'; 
signal C_4_S_1_L_0_out : std_logic := '0'; 
signal C_4_S_1_L_1_out : std_logic := '0'; 
signal C_4_S_1_L_2_out : std_logic := '0'; 
signal C_4_S_1_L_3_out : std_logic := '0'; 
signal C_4_S_1_L_4_out : std_logic := '0'; 
signal C_4_S_1_L_5_out : std_logic := '0'; 
signal C_4_S_1_L_6_out : std_logic := '0'; 
signal C_4_S_1_L_7_out : std_logic := '0'; 
signal C_4_S_2_L_0_out : std_logic := '0'; 
signal C_4_S_2_L_1_out : std_logic := '0'; 
signal C_4_S_2_L_2_out : std_logic := '0'; 
signal C_4_S_2_L_3_out : std_logic := '0'; 
signal C_4_S_2_L_4_out : std_logic := '0'; 
signal C_4_S_2_L_5_out : std_logic := '0'; 
signal C_4_S_2_L_6_out : std_logic := '0'; 
signal C_4_S_2_L_7_out : std_logic := '0'; 
signal C_4_S_3_L_0_out : std_logic := '0'; 
signal C_4_S_3_L_1_out : std_logic := '0'; 
signal C_4_S_3_L_2_out : std_logic := '0'; 
signal C_4_S_3_L_3_out : std_logic := '0'; 
signal C_4_S_3_L_4_out : std_logic := '0'; 
signal C_4_S_3_L_5_out : std_logic := '0'; 
signal C_4_S_3_L_6_out : std_logic := '0'; 
signal C_4_S_3_L_7_out : std_logic := '0'; 
signal C_4_S_4_L_0_out : std_logic := '0'; 
signal C_4_S_4_L_1_out : std_logic := '0'; 
signal C_4_S_4_L_2_out : std_logic := '0'; 
signal C_4_S_4_L_3_out : std_logic := '0'; 
signal C_4_S_4_L_4_out : std_logic := '0'; 
signal C_4_S_4_L_5_out : std_logic := '0'; 
signal C_4_S_4_L_6_out : std_logic := '0'; 
signal C_4_S_4_L_7_out : std_logic := '0'; 
signal C_5_S_0_L_0_out : std_logic := '0'; 
signal C_5_S_0_L_1_out : std_logic := '0'; 
signal C_5_S_0_L_2_out : std_logic := '0'; 
signal C_5_S_0_L_3_out : std_logic := '0'; 
signal C_5_S_0_L_4_out : std_logic := '0'; 
signal C_5_S_0_L_5_out : std_logic := '0'; 
signal C_5_S_0_L_6_out : std_logic := '0'; 
signal C_5_S_0_L_7_out : std_logic := '0'; 
signal C_5_S_1_L_0_out : std_logic := '0'; 
signal C_5_S_1_L_1_out : std_logic := '0'; 
signal C_5_S_1_L_2_out : std_logic := '0'; 
signal C_5_S_1_L_3_out : std_logic := '0'; 
signal C_5_S_1_L_4_out : std_logic := '0'; 
signal C_5_S_1_L_5_out : std_logic := '0'; 
signal C_5_S_1_L_6_out : std_logic := '0'; 
signal C_5_S_1_L_7_out : std_logic := '0'; 
signal C_5_S_2_L_0_out : std_logic := '0'; 
signal C_5_S_2_L_1_out : std_logic := '0'; 
signal C_5_S_2_L_2_out : std_logic := '0'; 
signal C_5_S_2_L_3_out : std_logic := '0'; 
signal C_5_S_2_L_4_out : std_logic := '0'; 
signal C_5_S_2_L_5_out : std_logic := '0'; 
signal C_5_S_2_L_6_out : std_logic := '0'; 
signal C_5_S_2_L_7_out : std_logic := '0'; 
signal C_5_S_3_L_0_out : std_logic := '0'; 
signal C_5_S_3_L_1_out : std_logic := '0'; 
signal C_5_S_3_L_2_out : std_logic := '0'; 
signal C_5_S_3_L_3_out : std_logic := '0'; 
signal C_5_S_3_L_4_out : std_logic := '0'; 
signal C_5_S_3_L_5_out : std_logic := '0'; 
signal C_5_S_3_L_6_out : std_logic := '0'; 
signal C_5_S_3_L_7_out : std_logic := '0'; 
signal C_5_S_4_L_0_out : std_logic := '0'; 
signal C_5_S_4_L_1_out : std_logic := '0'; 
signal C_5_S_4_L_2_out : std_logic := '0'; 
signal C_5_S_4_L_3_out : std_logic := '0'; 
signal C_5_S_4_L_4_out : std_logic := '0'; 
signal C_5_S_4_L_5_out : std_logic := '0'; 
signal C_5_S_4_L_6_out : std_logic := '0'; 
signal C_5_S_4_L_7_out : std_logic := '0'; 
signal C_6_S_0_L_0_out : std_logic := '0'; 
signal C_6_S_0_L_1_out : std_logic := '0'; 
signal C_6_S_0_L_2_out : std_logic := '0'; 
signal C_6_S_0_L_3_out : std_logic := '0'; 
signal C_6_S_0_L_4_out : std_logic := '0'; 
signal C_6_S_0_L_5_out : std_logic := '0'; 
signal C_6_S_0_L_6_out : std_logic := '0'; 
signal C_6_S_0_L_7_out : std_logic := '0'; 
signal C_6_S_1_L_0_out : std_logic := '0'; 
signal C_6_S_1_L_1_out : std_logic := '0'; 
signal C_6_S_1_L_2_out : std_logic := '0'; 
signal C_6_S_1_L_3_out : std_logic := '0'; 
signal C_6_S_1_L_4_out : std_logic := '0'; 
signal C_6_S_1_L_5_out : std_logic := '0'; 
signal C_6_S_1_L_6_out : std_logic := '0'; 
signal C_6_S_1_L_7_out : std_logic := '0'; 
signal C_6_S_2_L_0_out : std_logic := '0'; 
signal C_6_S_2_L_1_out : std_logic := '0'; 
signal C_6_S_2_L_2_out : std_logic := '0'; 
signal C_6_S_2_L_3_out : std_logic := '0'; 
signal C_6_S_2_L_4_out : std_logic := '0'; 
signal C_6_S_2_L_5_out : std_logic := '0'; 
signal C_6_S_2_L_6_out : std_logic := '0'; 
signal C_6_S_2_L_7_out : std_logic := '0'; 
signal C_6_S_3_L_0_out : std_logic := '0'; 
signal C_6_S_3_L_1_out : std_logic := '0'; 
signal C_6_S_3_L_2_out : std_logic := '0'; 
signal C_6_S_3_L_3_out : std_logic := '0'; 
signal C_6_S_3_L_4_out : std_logic := '0'; 
signal C_6_S_3_L_5_out : std_logic := '0'; 
signal C_6_S_3_L_6_out : std_logic := '0'; 
signal C_6_S_3_L_7_out : std_logic := '0'; 
signal C_6_S_4_L_0_out : std_logic := '0'; 
signal C_6_S_4_L_1_out : std_logic := '0'; 
signal C_6_S_4_L_2_out : std_logic := '0'; 
signal C_6_S_4_L_3_out : std_logic := '0'; 
signal C_6_S_4_L_4_out : std_logic := '0'; 
signal C_6_S_4_L_5_out : std_logic := '0'; 
signal C_6_S_4_L_6_out : std_logic := '0'; 
signal C_6_S_4_L_7_out : std_logic := '0'; 
signal C_7_S_0_L_0_out : std_logic := '0'; 
signal C_7_S_0_L_1_out : std_logic := '0'; 
signal C_7_S_0_L_2_out : std_logic := '0'; 
signal C_7_S_0_L_3_out : std_logic := '0'; 
signal C_7_S_0_L_4_out : std_logic := '0'; 
signal C_7_S_0_L_5_out : std_logic := '0'; 
signal C_7_S_0_L_6_out : std_logic := '0'; 
signal C_7_S_0_L_7_out : std_logic := '0'; 
signal C_7_S_1_L_0_out : std_logic := '0'; 
signal C_7_S_1_L_1_out : std_logic := '0'; 
signal C_7_S_1_L_2_out : std_logic := '0'; 
signal C_7_S_1_L_3_out : std_logic := '0'; 
signal C_7_S_1_L_4_out : std_logic := '0'; 
signal C_7_S_1_L_5_out : std_logic := '0'; 
signal C_7_S_1_L_6_out : std_logic := '0'; 
signal C_7_S_1_L_7_out : std_logic := '0'; 
signal C_7_S_2_L_0_out : std_logic := '0'; 
signal C_7_S_2_L_1_out : std_logic := '0'; 
signal C_7_S_2_L_2_out : std_logic := '0'; 
signal C_7_S_2_L_3_out : std_logic := '0'; 
signal C_7_S_2_L_4_out : std_logic := '0'; 
signal C_7_S_2_L_5_out : std_logic := '0'; 
signal C_7_S_2_L_6_out : std_logic := '0'; 
signal C_7_S_2_L_7_out : std_logic := '0'; 
signal C_7_S_3_L_0_out : std_logic := '0'; 
signal C_7_S_3_L_1_out : std_logic := '0'; 
signal C_7_S_3_L_2_out : std_logic := '0'; 
signal C_7_S_3_L_3_out : std_logic := '0'; 
signal C_7_S_3_L_4_out : std_logic := '0'; 
signal C_7_S_3_L_5_out : std_logic := '0'; 
signal C_7_S_3_L_6_out : std_logic := '0'; 
signal C_7_S_3_L_7_out : std_logic := '0'; 
signal C_7_S_4_L_0_out : std_logic := '0'; 
signal C_7_S_4_L_1_out : std_logic := '0'; 
signal C_7_S_4_L_2_out : std_logic := '0'; 
signal C_7_S_4_L_3_out : std_logic := '0'; 
signal C_7_S_4_L_4_out : std_logic := '0'; 
signal C_7_S_4_L_5_out : std_logic := '0'; 
signal C_7_S_4_L_6_out : std_logic := '0'; 
signal C_7_S_4_L_7_out : std_logic := '0'; 
signal C_8_S_0_L_0_out : std_logic := '0'; 
signal C_8_S_0_L_1_out : std_logic := '0'; 
signal C_8_S_0_L_2_out : std_logic := '0'; 
signal C_8_S_0_L_3_out : std_logic := '0'; 
signal C_8_S_0_L_4_out : std_logic := '0'; 
signal C_8_S_0_L_5_out : std_logic := '0'; 
signal C_8_S_0_L_6_out : std_logic := '0'; 
signal C_8_S_0_L_7_out : std_logic := '0'; 
signal C_8_S_1_L_0_out : std_logic := '0'; 
signal C_8_S_1_L_1_out : std_logic := '0'; 
signal C_8_S_1_L_2_out : std_logic := '0'; 
signal C_8_S_1_L_3_out : std_logic := '0'; 
signal C_8_S_1_L_4_out : std_logic := '0'; 
signal C_8_S_1_L_5_out : std_logic := '0'; 
signal C_8_S_1_L_6_out : std_logic := '0'; 
signal C_8_S_1_L_7_out : std_logic := '0'; 
signal C_8_S_2_L_0_out : std_logic := '0'; 
signal C_8_S_2_L_1_out : std_logic := '0'; 
signal C_8_S_2_L_2_out : std_logic := '0'; 
signal C_8_S_2_L_3_out : std_logic := '0'; 
signal C_8_S_2_L_4_out : std_logic := '0'; 
signal C_8_S_2_L_5_out : std_logic := '0'; 
signal C_8_S_2_L_6_out : std_logic := '0'; 
signal C_8_S_2_L_7_out : std_logic := '0'; 
signal C_8_S_3_L_0_out : std_logic := '0'; 
signal C_8_S_3_L_1_out : std_logic := '0'; 
signal C_8_S_3_L_2_out : std_logic := '0'; 
signal C_8_S_3_L_3_out : std_logic := '0'; 
signal C_8_S_3_L_4_out : std_logic := '0'; 
signal C_8_S_3_L_5_out : std_logic := '0'; 
signal C_8_S_3_L_6_out : std_logic := '0'; 
signal C_8_S_3_L_7_out : std_logic := '0'; 
signal C_8_S_4_L_0_out : std_logic := '0'; 
signal C_8_S_4_L_1_out : std_logic := '0'; 
signal C_8_S_4_L_2_out : std_logic := '0'; 
signal C_8_S_4_L_3_out : std_logic := '0'; 
signal C_8_S_4_L_4_out : std_logic := '0'; 
signal C_8_S_4_L_5_out : std_logic := '0'; 
signal C_8_S_4_L_6_out : std_logic := '0'; 
signal C_8_S_4_L_7_out : std_logic := '0'; 
signal C_9_S_0_L_0_out : std_logic := '0'; 
signal C_9_S_0_L_1_out : std_logic := '0'; 
signal C_9_S_0_L_2_out : std_logic := '0'; 
signal C_9_S_0_L_3_out : std_logic := '0'; 
signal C_9_S_0_L_4_out : std_logic := '0'; 
signal C_9_S_0_L_5_out : std_logic := '0'; 
signal C_9_S_0_L_6_out : std_logic := '0'; 
signal C_9_S_0_L_7_out : std_logic := '0'; 
signal C_9_S_1_L_0_out : std_logic := '0'; 
signal C_9_S_1_L_1_out : std_logic := '0'; 
signal C_9_S_1_L_2_out : std_logic := '0'; 
signal C_9_S_1_L_3_out : std_logic := '0'; 
signal C_9_S_1_L_4_out : std_logic := '0'; 
signal C_9_S_1_L_5_out : std_logic := '0'; 
signal C_9_S_1_L_6_out : std_logic := '0'; 
signal C_9_S_1_L_7_out : std_logic := '0'; 
signal C_9_S_2_L_0_out : std_logic := '0'; 
signal C_9_S_2_L_1_out : std_logic := '0'; 
signal C_9_S_2_L_2_out : std_logic := '0'; 
signal C_9_S_2_L_3_out : std_logic := '0'; 
signal C_9_S_2_L_4_out : std_logic := '0'; 
signal C_9_S_2_L_5_out : std_logic := '0'; 
signal C_9_S_2_L_6_out : std_logic := '0'; 
signal C_9_S_2_L_7_out : std_logic := '0'; 
signal C_9_S_3_L_0_out : std_logic := '0'; 
signal C_9_S_3_L_1_out : std_logic := '0'; 
signal C_9_S_3_L_2_out : std_logic := '0'; 
signal C_9_S_3_L_3_out : std_logic := '0'; 
signal C_9_S_3_L_4_out : std_logic := '0'; 
signal C_9_S_3_L_5_out : std_logic := '0'; 
signal C_9_S_3_L_6_out : std_logic := '0'; 
signal C_9_S_3_L_7_out : std_logic := '0'; 
signal C_9_S_4_L_0_out : std_logic := '0'; 
signal C_9_S_4_L_1_out : std_logic := '0'; 
signal C_9_S_4_L_2_out : std_logic := '0'; 
signal C_9_S_4_L_3_out : std_logic := '0'; 
signal C_9_S_4_L_4_out : std_logic := '0'; 
signal C_9_S_4_L_5_out : std_logic := '0'; 
signal C_9_S_4_L_6_out : std_logic := '0'; 
signal C_9_S_4_L_7_out : std_logic := '0'; 
signal C_10_S_0_L_0_out : std_logic := '0'; 
signal C_10_S_0_L_1_out : std_logic := '0'; 
signal C_10_S_0_L_2_out : std_logic := '0'; 
signal C_10_S_0_L_3_out : std_logic := '0'; 
signal C_10_S_0_L_4_out : std_logic := '0'; 
signal C_10_S_0_L_5_out : std_logic := '0'; 
signal C_10_S_0_L_6_out : std_logic := '0'; 
signal C_10_S_0_L_7_out : std_logic := '0'; 
signal C_10_S_1_L_0_out : std_logic := '0'; 
signal C_10_S_1_L_1_out : std_logic := '0'; 
signal C_10_S_1_L_2_out : std_logic := '0'; 
signal C_10_S_1_L_3_out : std_logic := '0'; 
signal C_10_S_1_L_4_out : std_logic := '0'; 
signal C_10_S_1_L_5_out : std_logic := '0'; 
signal C_10_S_1_L_6_out : std_logic := '0'; 
signal C_10_S_1_L_7_out : std_logic := '0'; 
signal C_10_S_2_L_0_out : std_logic := '0'; 
signal C_10_S_2_L_1_out : std_logic := '0'; 
signal C_10_S_2_L_2_out : std_logic := '0'; 
signal C_10_S_2_L_3_out : std_logic := '0'; 
signal C_10_S_2_L_4_out : std_logic := '0'; 
signal C_10_S_2_L_5_out : std_logic := '0'; 
signal C_10_S_2_L_6_out : std_logic := '0'; 
signal C_10_S_2_L_7_out : std_logic := '0'; 
signal C_10_S_3_L_0_out : std_logic := '0'; 
signal C_10_S_3_L_1_out : std_logic := '0'; 
signal C_10_S_3_L_2_out : std_logic := '0'; 
signal C_10_S_3_L_3_out : std_logic := '0'; 
signal C_10_S_3_L_4_out : std_logic := '0'; 
signal C_10_S_3_L_5_out : std_logic := '0'; 
signal C_10_S_3_L_6_out : std_logic := '0'; 
signal C_10_S_3_L_7_out : std_logic := '0'; 
signal C_10_S_4_L_0_out : std_logic := '0'; 
signal C_10_S_4_L_1_out : std_logic := '0'; 
signal C_10_S_4_L_2_out : std_logic := '0'; 
signal C_10_S_4_L_3_out : std_logic := '0'; 
signal C_10_S_4_L_4_out : std_logic := '0'; 
signal C_10_S_4_L_5_out : std_logic := '0'; 
signal C_10_S_4_L_6_out : std_logic := '0'; 
signal C_10_S_4_L_7_out : std_logic := '0'; 
signal C_11_S_0_L_0_out : std_logic := '0'; 
signal C_11_S_0_L_1_out : std_logic := '0'; 
signal C_11_S_0_L_2_out : std_logic := '0'; 
signal C_11_S_0_L_3_out : std_logic := '0'; 
signal C_11_S_0_L_4_out : std_logic := '0'; 
signal C_11_S_0_L_5_out : std_logic := '0'; 
signal C_11_S_0_L_6_out : std_logic := '0'; 
signal C_11_S_0_L_7_out : std_logic := '0'; 
signal C_11_S_1_L_0_out : std_logic := '0'; 
signal C_11_S_1_L_1_out : std_logic := '0'; 
signal C_11_S_1_L_2_out : std_logic := '0'; 
signal C_11_S_1_L_3_out : std_logic := '0'; 
signal C_11_S_1_L_4_out : std_logic := '0'; 
signal C_11_S_1_L_5_out : std_logic := '0'; 
signal C_11_S_1_L_6_out : std_logic := '0'; 
signal C_11_S_1_L_7_out : std_logic := '0'; 
signal C_11_S_2_L_0_out : std_logic := '0'; 
signal C_11_S_2_L_1_out : std_logic := '0'; 
signal C_11_S_2_L_2_out : std_logic := '0'; 
signal C_11_S_2_L_3_out : std_logic := '0'; 
signal C_11_S_2_L_4_out : std_logic := '0'; 
signal C_11_S_2_L_5_out : std_logic := '0'; 
signal C_11_S_2_L_6_out : std_logic := '0'; 
signal C_11_S_2_L_7_out : std_logic := '0'; 
signal C_11_S_3_L_0_out : std_logic := '0'; 
signal C_11_S_3_L_1_out : std_logic := '0'; 
signal C_11_S_3_L_2_out : std_logic := '0'; 
signal C_11_S_3_L_3_out : std_logic := '0'; 
signal C_11_S_3_L_4_out : std_logic := '0'; 
signal C_11_S_3_L_5_out : std_logic := '0'; 
signal C_11_S_3_L_6_out : std_logic := '0'; 
signal C_11_S_3_L_7_out : std_logic := '0'; 
signal C_11_S_4_L_0_out : std_logic := '0'; 
signal C_11_S_4_L_1_out : std_logic := '0'; 
signal C_11_S_4_L_2_out : std_logic := '0'; 
signal C_11_S_4_L_3_out : std_logic := '0'; 
signal C_11_S_4_L_4_out : std_logic := '0'; 
signal C_11_S_4_L_5_out : std_logic := '0'; 
signal C_11_S_4_L_6_out : std_logic := '0'; 
signal C_11_S_4_L_7_out : std_logic := '0'; 
signal C_12_S_0_L_0_out : std_logic := '0'; 
signal C_12_S_0_L_1_out : std_logic := '0'; 
signal C_12_S_0_L_2_out : std_logic := '0'; 
signal C_12_S_0_L_3_out : std_logic := '0'; 
signal C_12_S_0_L_4_out : std_logic := '0'; 
signal C_12_S_0_L_5_out : std_logic := '0'; 
signal C_12_S_0_L_6_out : std_logic := '0'; 
signal C_12_S_0_L_7_out : std_logic := '0'; 
signal C_12_S_1_L_0_out : std_logic := '0'; 
signal C_12_S_1_L_1_out : std_logic := '0'; 
signal C_12_S_1_L_2_out : std_logic := '0'; 
signal C_12_S_1_L_3_out : std_logic := '0'; 
signal C_12_S_1_L_4_out : std_logic := '0'; 
signal C_12_S_1_L_5_out : std_logic := '0'; 
signal C_12_S_1_L_6_out : std_logic := '0'; 
signal C_12_S_1_L_7_out : std_logic := '0'; 
signal C_12_S_2_L_0_out : std_logic := '0'; 
signal C_12_S_2_L_1_out : std_logic := '0'; 
signal C_12_S_2_L_2_out : std_logic := '0'; 
signal C_12_S_2_L_3_out : std_logic := '0'; 
signal C_12_S_2_L_4_out : std_logic := '0'; 
signal C_12_S_2_L_5_out : std_logic := '0'; 
signal C_12_S_2_L_6_out : std_logic := '0'; 
signal C_12_S_2_L_7_out : std_logic := '0'; 
signal C_12_S_3_L_0_out : std_logic := '0'; 
signal C_12_S_3_L_1_out : std_logic := '0'; 
signal C_12_S_3_L_2_out : std_logic := '0'; 
signal C_12_S_3_L_3_out : std_logic := '0'; 
signal C_12_S_3_L_4_out : std_logic := '0'; 
signal C_12_S_3_L_5_out : std_logic := '0'; 
signal C_12_S_3_L_6_out : std_logic := '0'; 
signal C_12_S_3_L_7_out : std_logic := '0'; 
signal C_12_S_4_L_0_out : std_logic := '0'; 
signal C_12_S_4_L_1_out : std_logic := '0'; 
signal C_12_S_4_L_2_out : std_logic := '0'; 
signal C_12_S_4_L_3_out : std_logic := '0'; 
signal C_12_S_4_L_4_out : std_logic := '0'; 
signal C_12_S_4_L_5_out : std_logic := '0'; 
signal C_12_S_4_L_6_out : std_logic := '0'; 
signal C_12_S_4_L_7_out : std_logic := '0'; 
signal C_13_S_0_L_0_out : std_logic := '0'; 
signal C_13_S_0_L_1_out : std_logic := '0'; 
signal C_13_S_0_L_2_out : std_logic := '0'; 
signal C_13_S_0_L_3_out : std_logic := '0'; 
signal C_13_S_0_L_4_out : std_logic := '0'; 
signal C_13_S_0_L_5_out : std_logic := '0'; 
signal C_13_S_0_L_6_out : std_logic := '0'; 
signal C_13_S_0_L_7_out : std_logic := '0'; 
signal C_13_S_1_L_0_out : std_logic := '0'; 
signal C_13_S_1_L_1_out : std_logic := '0'; 
signal C_13_S_1_L_2_out : std_logic := '0'; 
signal C_13_S_1_L_3_out : std_logic := '0'; 
signal C_13_S_1_L_4_out : std_logic := '0'; 
signal C_13_S_1_L_5_out : std_logic := '0'; 
signal C_13_S_1_L_6_out : std_logic := '0'; 
signal C_13_S_1_L_7_out : std_logic := '0'; 
signal C_13_S_2_L_0_out : std_logic := '0'; 
signal C_13_S_2_L_1_out : std_logic := '0'; 
signal C_13_S_2_L_2_out : std_logic := '0'; 
signal C_13_S_2_L_3_out : std_logic := '0'; 
signal C_13_S_2_L_4_out : std_logic := '0'; 
signal C_13_S_2_L_5_out : std_logic := '0'; 
signal C_13_S_2_L_6_out : std_logic := '0'; 
signal C_13_S_2_L_7_out : std_logic := '0'; 
signal C_13_S_3_L_0_out : std_logic := '0'; 
signal C_13_S_3_L_1_out : std_logic := '0'; 
signal C_13_S_3_L_2_out : std_logic := '0'; 
signal C_13_S_3_L_3_out : std_logic := '0'; 
signal C_13_S_3_L_4_out : std_logic := '0'; 
signal C_13_S_3_L_5_out : std_logic := '0'; 
signal C_13_S_3_L_6_out : std_logic := '0'; 
signal C_13_S_3_L_7_out : std_logic := '0'; 
signal C_13_S_4_L_0_out : std_logic := '0'; 
signal C_13_S_4_L_1_out : std_logic := '0'; 
signal C_13_S_4_L_2_out : std_logic := '0'; 
signal C_13_S_4_L_3_out : std_logic := '0'; 
signal C_13_S_4_L_4_out : std_logic := '0'; 
signal C_13_S_4_L_5_out : std_logic := '0'; 
signal C_13_S_4_L_6_out : std_logic := '0'; 
signal C_13_S_4_L_7_out : std_logic := '0'; 
signal C_14_S_0_L_0_out : std_logic := '0'; 
signal C_14_S_0_L_1_out : std_logic := '0'; 
signal C_14_S_0_L_2_out : std_logic := '0'; 
signal C_14_S_0_L_3_out : std_logic := '0'; 
signal C_14_S_0_L_4_out : std_logic := '0'; 
signal C_14_S_0_L_5_out : std_logic := '0'; 
signal C_14_S_0_L_6_out : std_logic := '0'; 
signal C_14_S_0_L_7_out : std_logic := '0'; 
signal C_14_S_1_L_0_out : std_logic := '0'; 
signal C_14_S_1_L_1_out : std_logic := '0'; 
signal C_14_S_1_L_2_out : std_logic := '0'; 
signal C_14_S_1_L_3_out : std_logic := '0'; 
signal C_14_S_1_L_4_out : std_logic := '0'; 
signal C_14_S_1_L_5_out : std_logic := '0'; 
signal C_14_S_1_L_6_out : std_logic := '0'; 
signal C_14_S_1_L_7_out : std_logic := '0'; 
signal C_14_S_2_L_0_out : std_logic := '0'; 
signal C_14_S_2_L_1_out : std_logic := '0'; 
signal C_14_S_2_L_2_out : std_logic := '0'; 
signal C_14_S_2_L_3_out : std_logic := '0'; 
signal C_14_S_2_L_4_out : std_logic := '0'; 
signal C_14_S_2_L_5_out : std_logic := '0'; 
signal C_14_S_2_L_6_out : std_logic := '0'; 
signal C_14_S_2_L_7_out : std_logic := '0'; 
signal C_14_S_3_L_0_out : std_logic := '0'; 
signal C_14_S_3_L_1_out : std_logic := '0'; 
signal C_14_S_3_L_2_out : std_logic := '0'; 
signal C_14_S_3_L_3_out : std_logic := '0'; 
signal C_14_S_3_L_4_out : std_logic := '0'; 
signal C_14_S_3_L_5_out : std_logic := '0'; 
signal C_14_S_3_L_6_out : std_logic := '0'; 
signal C_14_S_3_L_7_out : std_logic := '0'; 
signal C_14_S_4_L_0_out : std_logic := '0'; 
signal C_14_S_4_L_1_out : std_logic := '0'; 
signal C_14_S_4_L_2_out : std_logic := '0'; 
signal C_14_S_4_L_3_out : std_logic := '0'; 
signal C_14_S_4_L_4_out : std_logic := '0'; 
signal C_14_S_4_L_5_out : std_logic := '0'; 
signal C_14_S_4_L_6_out : std_logic := '0'; 
signal C_14_S_4_L_7_out : std_logic := '0'; 
signal C_15_S_0_L_0_out : std_logic := '0'; 
signal C_15_S_0_L_1_out : std_logic := '0'; 
signal C_15_S_0_L_2_out : std_logic := '0'; 
signal C_15_S_0_L_3_out : std_logic := '0'; 
signal C_15_S_0_L_4_out : std_logic := '0'; 
signal C_15_S_0_L_5_out : std_logic := '0'; 
signal C_15_S_0_L_6_out : std_logic := '0'; 
signal C_15_S_0_L_7_out : std_logic := '0'; 
signal C_15_S_1_L_0_out : std_logic := '0'; 
signal C_15_S_1_L_1_out : std_logic := '0'; 
signal C_15_S_1_L_2_out : std_logic := '0'; 
signal C_15_S_1_L_3_out : std_logic := '0'; 
signal C_15_S_1_L_4_out : std_logic := '0'; 
signal C_15_S_1_L_5_out : std_logic := '0'; 
signal C_15_S_1_L_6_out : std_logic := '0'; 
signal C_15_S_1_L_7_out : std_logic := '0'; 
signal C_15_S_2_L_0_out : std_logic := '0'; 
signal C_15_S_2_L_1_out : std_logic := '0'; 
signal C_15_S_2_L_2_out : std_logic := '0'; 
signal C_15_S_2_L_3_out : std_logic := '0'; 
signal C_15_S_2_L_4_out : std_logic := '0'; 
signal C_15_S_2_L_5_out : std_logic := '0'; 
signal C_15_S_2_L_6_out : std_logic := '0'; 
signal C_15_S_2_L_7_out : std_logic := '0'; 
signal C_15_S_3_L_0_out : std_logic := '0'; 
signal C_15_S_3_L_1_out : std_logic := '0'; 
signal C_15_S_3_L_2_out : std_logic := '0'; 
signal C_15_S_3_L_3_out : std_logic := '0'; 
signal C_15_S_3_L_4_out : std_logic := '0'; 
signal C_15_S_3_L_5_out : std_logic := '0'; 
signal C_15_S_3_L_6_out : std_logic := '0'; 
signal C_15_S_3_L_7_out : std_logic := '0'; 
signal C_15_S_4_L_0_out : std_logic := '0'; 
signal C_15_S_4_L_1_out : std_logic := '0'; 
signal C_15_S_4_L_2_out : std_logic := '0'; 
signal C_15_S_4_L_3_out : std_logic := '0'; 
signal C_15_S_4_L_4_out : std_logic := '0'; 
signal C_15_S_4_L_5_out : std_logic := '0'; 
signal C_15_S_4_L_6_out : std_logic := '0'; 
signal C_15_S_4_L_7_out : std_logic := '0'; 
signal C_16_S_0_L_0_out : std_logic := '0'; 
signal C_16_S_0_L_1_out : std_logic := '0'; 
signal C_16_S_0_L_2_out : std_logic := '0'; 
signal C_16_S_0_L_3_out : std_logic := '0'; 
signal C_16_S_0_L_4_out : std_logic := '0'; 
signal C_16_S_0_L_5_out : std_logic := '0'; 
signal C_16_S_0_L_6_out : std_logic := '0'; 
signal C_16_S_0_L_7_out : std_logic := '0'; 
signal C_16_S_1_L_0_out : std_logic := '0'; 
signal C_16_S_1_L_1_out : std_logic := '0'; 
signal C_16_S_1_L_2_out : std_logic := '0'; 
signal C_16_S_1_L_3_out : std_logic := '0'; 
signal C_16_S_1_L_4_out : std_logic := '0'; 
signal C_16_S_1_L_5_out : std_logic := '0'; 
signal C_16_S_1_L_6_out : std_logic := '0'; 
signal C_16_S_1_L_7_out : std_logic := '0'; 
signal C_16_S_2_L_0_out : std_logic := '0'; 
signal C_16_S_2_L_1_out : std_logic := '0'; 
signal C_16_S_2_L_2_out : std_logic := '0'; 
signal C_16_S_2_L_3_out : std_logic := '0'; 
signal C_16_S_2_L_4_out : std_logic := '0'; 
signal C_16_S_2_L_5_out : std_logic := '0'; 
signal C_16_S_2_L_6_out : std_logic := '0'; 
signal C_16_S_2_L_7_out : std_logic := '0'; 
signal C_16_S_3_L_0_out : std_logic := '0'; 
signal C_16_S_3_L_1_out : std_logic := '0'; 
signal C_16_S_3_L_2_out : std_logic := '0'; 
signal C_16_S_3_L_3_out : std_logic := '0'; 
signal C_16_S_3_L_4_out : std_logic := '0'; 
signal C_16_S_3_L_5_out : std_logic := '0'; 
signal C_16_S_3_L_6_out : std_logic := '0'; 
signal C_16_S_3_L_7_out : std_logic := '0'; 
signal C_16_S_4_L_0_out : std_logic := '0'; 
signal C_16_S_4_L_1_out : std_logic := '0'; 
signal C_16_S_4_L_2_out : std_logic := '0'; 
signal C_16_S_4_L_3_out : std_logic := '0'; 
signal C_16_S_4_L_4_out : std_logic := '0'; 
signal C_16_S_4_L_5_out : std_logic := '0'; 
signal C_16_S_4_L_6_out : std_logic := '0'; 
signal C_16_S_4_L_7_out : std_logic := '0'; 
signal C_17_S_0_L_0_out : std_logic := '0'; 
signal C_17_S_0_L_1_out : std_logic := '0'; 
signal C_17_S_0_L_2_out : std_logic := '0'; 
signal C_17_S_0_L_3_out : std_logic := '0'; 
signal C_17_S_0_L_4_out : std_logic := '0'; 
signal C_17_S_0_L_5_out : std_logic := '0'; 
signal C_17_S_0_L_6_out : std_logic := '0'; 
signal C_17_S_0_L_7_out : std_logic := '0'; 
signal C_17_S_1_L_0_out : std_logic := '0'; 
signal C_17_S_1_L_1_out : std_logic := '0'; 
signal C_17_S_1_L_2_out : std_logic := '0'; 
signal C_17_S_1_L_3_out : std_logic := '0'; 
signal C_17_S_1_L_4_out : std_logic := '0'; 
signal C_17_S_1_L_5_out : std_logic := '0'; 
signal C_17_S_1_L_6_out : std_logic := '0'; 
signal C_17_S_1_L_7_out : std_logic := '0'; 
signal C_17_S_2_L_0_out : std_logic := '0'; 
signal C_17_S_2_L_1_out : std_logic := '0'; 
signal C_17_S_2_L_2_out : std_logic := '0'; 
signal C_17_S_2_L_3_out : std_logic := '0'; 
signal C_17_S_2_L_4_out : std_logic := '0'; 
signal C_17_S_2_L_5_out : std_logic := '0'; 
signal C_17_S_2_L_6_out : std_logic := '0'; 
signal C_17_S_2_L_7_out : std_logic := '0'; 
signal C_17_S_3_L_0_out : std_logic := '0'; 
signal C_17_S_3_L_1_out : std_logic := '0'; 
signal C_17_S_3_L_2_out : std_logic := '0'; 
signal C_17_S_3_L_3_out : std_logic := '0'; 
signal C_17_S_3_L_4_out : std_logic := '0'; 
signal C_17_S_3_L_5_out : std_logic := '0'; 
signal C_17_S_3_L_6_out : std_logic := '0'; 
signal C_17_S_3_L_7_out : std_logic := '0'; 
signal C_17_S_4_L_0_out : std_logic := '0'; 
signal C_17_S_4_L_1_out : std_logic := '0'; 
signal C_17_S_4_L_2_out : std_logic := '0'; 
signal C_17_S_4_L_3_out : std_logic := '0'; 
signal C_17_S_4_L_4_out : std_logic := '0'; 
signal C_17_S_4_L_5_out : std_logic := '0'; 
signal C_17_S_4_L_6_out : std_logic := '0'; 
signal C_17_S_4_L_7_out : std_logic := '0'; 
signal C_18_S_0_L_0_out : std_logic := '0'; 
signal C_18_S_0_L_1_out : std_logic := '0'; 
signal C_18_S_0_L_2_out : std_logic := '0'; 
signal C_18_S_0_L_3_out : std_logic := '0'; 
signal C_18_S_0_L_4_out : std_logic := '0'; 
signal C_18_S_0_L_5_out : std_logic := '0'; 
signal C_18_S_0_L_6_out : std_logic := '0'; 
signal C_18_S_0_L_7_out : std_logic := '0'; 
signal C_18_S_1_L_0_out : std_logic := '0'; 
signal C_18_S_1_L_1_out : std_logic := '0'; 
signal C_18_S_1_L_2_out : std_logic := '0'; 
signal C_18_S_1_L_3_out : std_logic := '0'; 
signal C_18_S_1_L_4_out : std_logic := '0'; 
signal C_18_S_1_L_5_out : std_logic := '0'; 
signal C_18_S_1_L_6_out : std_logic := '0'; 
signal C_18_S_1_L_7_out : std_logic := '0'; 
signal C_18_S_2_L_0_out : std_logic := '0'; 
signal C_18_S_2_L_1_out : std_logic := '0'; 
signal C_18_S_2_L_2_out : std_logic := '0'; 
signal C_18_S_2_L_3_out : std_logic := '0'; 
signal C_18_S_2_L_4_out : std_logic := '0'; 
signal C_18_S_2_L_5_out : std_logic := '0'; 
signal C_18_S_2_L_6_out : std_logic := '0'; 
signal C_18_S_2_L_7_out : std_logic := '0'; 
signal C_18_S_3_L_0_out : std_logic := '0'; 
signal C_18_S_3_L_1_out : std_logic := '0'; 
signal C_18_S_3_L_2_out : std_logic := '0'; 
signal C_18_S_3_L_3_out : std_logic := '0'; 
signal C_18_S_3_L_4_out : std_logic := '0'; 
signal C_18_S_3_L_5_out : std_logic := '0'; 
signal C_18_S_3_L_6_out : std_logic := '0'; 
signal C_18_S_3_L_7_out : std_logic := '0'; 
signal C_18_S_4_L_0_out : std_logic := '0'; 
signal C_18_S_4_L_1_out : std_logic := '0'; 
signal C_18_S_4_L_2_out : std_logic := '0'; 
signal C_18_S_4_L_3_out : std_logic := '0'; 
signal C_18_S_4_L_4_out : std_logic := '0'; 
signal C_18_S_4_L_5_out : std_logic := '0'; 
signal C_18_S_4_L_6_out : std_logic := '0'; 
signal C_18_S_4_L_7_out : std_logic := '0'; 
signal C_19_S_0_L_0_out : std_logic := '0'; 
signal C_19_S_0_L_1_out : std_logic := '0'; 
signal C_19_S_0_L_2_out : std_logic := '0'; 
signal C_19_S_0_L_3_out : std_logic := '0'; 
signal C_19_S_0_L_4_out : std_logic := '0'; 
signal C_19_S_0_L_5_out : std_logic := '0'; 
signal C_19_S_0_L_6_out : std_logic := '0'; 
signal C_19_S_0_L_7_out : std_logic := '0'; 
signal C_19_S_1_L_0_out : std_logic := '0'; 
signal C_19_S_1_L_1_out : std_logic := '0'; 
signal C_19_S_1_L_2_out : std_logic := '0'; 
signal C_19_S_1_L_3_out : std_logic := '0'; 
signal C_19_S_1_L_4_out : std_logic := '0'; 
signal C_19_S_1_L_5_out : std_logic := '0'; 
signal C_19_S_1_L_6_out : std_logic := '0'; 
signal C_19_S_1_L_7_out : std_logic := '0'; 
signal C_19_S_2_L_0_out : std_logic := '0'; 
signal C_19_S_2_L_1_out : std_logic := '0'; 
signal C_19_S_2_L_2_out : std_logic := '0'; 
signal C_19_S_2_L_3_out : std_logic := '0'; 
signal C_19_S_2_L_4_out : std_logic := '0'; 
signal C_19_S_2_L_5_out : std_logic := '0'; 
signal C_19_S_2_L_6_out : std_logic := '0'; 
signal C_19_S_2_L_7_out : std_logic := '0'; 
signal C_19_S_3_L_0_out : std_logic := '0'; 
signal C_19_S_3_L_1_out : std_logic := '0'; 
signal C_19_S_3_L_2_out : std_logic := '0'; 
signal C_19_S_3_L_3_out : std_logic := '0'; 
signal C_19_S_3_L_4_out : std_logic := '0'; 
signal C_19_S_3_L_5_out : std_logic := '0'; 
signal C_19_S_3_L_6_out : std_logic := '0'; 
signal C_19_S_3_L_7_out : std_logic := '0'; 
signal C_19_S_4_L_0_out : std_logic := '0'; 
signal C_19_S_4_L_1_out : std_logic := '0'; 
signal C_19_S_4_L_2_out : std_logic := '0'; 
signal C_19_S_4_L_3_out : std_logic := '0'; 
signal C_19_S_4_L_4_out : std_logic := '0'; 
signal C_19_S_4_L_5_out : std_logic := '0'; 
signal C_19_S_4_L_6_out : std_logic := '0'; 
signal C_19_S_4_L_7_out : std_logic := '0'; 
signal C_20_S_0_L_0_out : std_logic := '0'; 
signal C_20_S_0_L_1_out : std_logic := '0'; 
signal C_20_S_0_L_2_out : std_logic := '0'; 
signal C_20_S_0_L_3_out : std_logic := '0'; 
signal C_20_S_0_L_4_out : std_logic := '0'; 
signal C_20_S_0_L_5_out : std_logic := '0'; 
signal C_20_S_0_L_6_out : std_logic := '0'; 
signal C_20_S_0_L_7_out : std_logic := '0'; 
signal C_20_S_1_L_0_out : std_logic := '0'; 
signal C_20_S_1_L_1_out : std_logic := '0'; 
signal C_20_S_1_L_2_out : std_logic := '0'; 
signal C_20_S_1_L_3_out : std_logic := '0'; 
signal C_20_S_1_L_4_out : std_logic := '0'; 
signal C_20_S_1_L_5_out : std_logic := '0'; 
signal C_20_S_1_L_6_out : std_logic := '0'; 
signal C_20_S_1_L_7_out : std_logic := '0'; 
signal C_20_S_2_L_0_out : std_logic := '0'; 
signal C_20_S_2_L_1_out : std_logic := '0'; 
signal C_20_S_2_L_2_out : std_logic := '0'; 
signal C_20_S_2_L_3_out : std_logic := '0'; 
signal C_20_S_2_L_4_out : std_logic := '0'; 
signal C_20_S_2_L_5_out : std_logic := '0'; 
signal C_20_S_2_L_6_out : std_logic := '0'; 
signal C_20_S_2_L_7_out : std_logic := '0'; 
signal C_20_S_3_L_0_out : std_logic := '0'; 
signal C_20_S_3_L_1_out : std_logic := '0'; 
signal C_20_S_3_L_2_out : std_logic := '0'; 
signal C_20_S_3_L_3_out : std_logic := '0'; 
signal C_20_S_3_L_4_out : std_logic := '0'; 
signal C_20_S_3_L_5_out : std_logic := '0'; 
signal C_20_S_3_L_6_out : std_logic := '0'; 
signal C_20_S_3_L_7_out : std_logic := '0'; 
signal C_20_S_4_L_0_out : std_logic := '0'; 
signal C_20_S_4_L_1_out : std_logic := '0'; 
signal C_20_S_4_L_2_out : std_logic := '0'; 
signal C_20_S_4_L_3_out : std_logic := '0'; 
signal C_20_S_4_L_4_out : std_logic := '0'; 
signal C_20_S_4_L_5_out : std_logic := '0'; 
signal C_20_S_4_L_6_out : std_logic := '0'; 
signal C_20_S_4_L_7_out : std_logic := '0'; 
signal C_21_S_0_L_0_out : std_logic := '0'; 
signal C_21_S_0_L_1_out : std_logic := '0'; 
signal C_21_S_0_L_2_out : std_logic := '0'; 
signal C_21_S_0_L_3_out : std_logic := '0'; 
signal C_21_S_0_L_4_out : std_logic := '0'; 
signal C_21_S_0_L_5_out : std_logic := '0'; 
signal C_21_S_0_L_6_out : std_logic := '0'; 
signal C_21_S_0_L_7_out : std_logic := '0'; 
signal C_21_S_1_L_0_out : std_logic := '0'; 
signal C_21_S_1_L_1_out : std_logic := '0'; 
signal C_21_S_1_L_2_out : std_logic := '0'; 
signal C_21_S_1_L_3_out : std_logic := '0'; 
signal C_21_S_1_L_4_out : std_logic := '0'; 
signal C_21_S_1_L_5_out : std_logic := '0'; 
signal C_21_S_1_L_6_out : std_logic := '0'; 
signal C_21_S_1_L_7_out : std_logic := '0'; 
signal C_21_S_2_L_0_out : std_logic := '0'; 
signal C_21_S_2_L_1_out : std_logic := '0'; 
signal C_21_S_2_L_2_out : std_logic := '0'; 
signal C_21_S_2_L_3_out : std_logic := '0'; 
signal C_21_S_2_L_4_out : std_logic := '0'; 
signal C_21_S_2_L_5_out : std_logic := '0'; 
signal C_21_S_2_L_6_out : std_logic := '0'; 
signal C_21_S_2_L_7_out : std_logic := '0'; 
signal C_21_S_3_L_0_out : std_logic := '0'; 
signal C_21_S_3_L_1_out : std_logic := '0'; 
signal C_21_S_3_L_2_out : std_logic := '0'; 
signal C_21_S_3_L_3_out : std_logic := '0'; 
signal C_21_S_3_L_4_out : std_logic := '0'; 
signal C_21_S_3_L_5_out : std_logic := '0'; 
signal C_21_S_3_L_6_out : std_logic := '0'; 
signal C_21_S_3_L_7_out : std_logic := '0'; 
signal C_21_S_4_L_0_out : std_logic := '0'; 
signal C_21_S_4_L_1_out : std_logic := '0'; 
signal C_21_S_4_L_2_out : std_logic := '0'; 
signal C_21_S_4_L_3_out : std_logic := '0'; 
signal C_21_S_4_L_4_out : std_logic := '0'; 
signal C_21_S_4_L_5_out : std_logic := '0'; 
signal C_21_S_4_L_6_out : std_logic := '0'; 
signal C_21_S_4_L_7_out : std_logic := '0'; 
signal C_22_S_0_L_0_out : std_logic := '0'; 
signal C_22_S_0_L_1_out : std_logic := '0'; 
signal C_22_S_0_L_2_out : std_logic := '0'; 
signal C_22_S_0_L_3_out : std_logic := '0'; 
signal C_22_S_0_L_4_out : std_logic := '0'; 
signal C_22_S_0_L_5_out : std_logic := '0'; 
signal C_22_S_0_L_6_out : std_logic := '0'; 
signal C_22_S_0_L_7_out : std_logic := '0'; 
signal C_22_S_1_L_0_out : std_logic := '0'; 
signal C_22_S_1_L_1_out : std_logic := '0'; 
signal C_22_S_1_L_2_out : std_logic := '0'; 
signal C_22_S_1_L_3_out : std_logic := '0'; 
signal C_22_S_1_L_4_out : std_logic := '0'; 
signal C_22_S_1_L_5_out : std_logic := '0'; 
signal C_22_S_1_L_6_out : std_logic := '0'; 
signal C_22_S_1_L_7_out : std_logic := '0'; 
signal C_22_S_2_L_0_out : std_logic := '0'; 
signal C_22_S_2_L_1_out : std_logic := '0'; 
signal C_22_S_2_L_2_out : std_logic := '0'; 
signal C_22_S_2_L_3_out : std_logic := '0'; 
signal C_22_S_2_L_4_out : std_logic := '0'; 
signal C_22_S_2_L_5_out : std_logic := '0'; 
signal C_22_S_2_L_6_out : std_logic := '0'; 
signal C_22_S_2_L_7_out : std_logic := '0'; 
signal C_22_S_3_L_0_out : std_logic := '0'; 
signal C_22_S_3_L_1_out : std_logic := '0'; 
signal C_22_S_3_L_2_out : std_logic := '0'; 
signal C_22_S_3_L_3_out : std_logic := '0'; 
signal C_22_S_3_L_4_out : std_logic := '0'; 
signal C_22_S_3_L_5_out : std_logic := '0'; 
signal C_22_S_3_L_6_out : std_logic := '0'; 
signal C_22_S_3_L_7_out : std_logic := '0'; 
signal C_22_S_4_L_0_out : std_logic := '0'; 
signal C_22_S_4_L_1_out : std_logic := '0'; 
signal C_22_S_4_L_2_out : std_logic := '0'; 
signal C_22_S_4_L_3_out : std_logic := '0'; 
signal C_22_S_4_L_4_out : std_logic := '0'; 
signal C_22_S_4_L_5_out : std_logic := '0'; 
signal C_22_S_4_L_6_out : std_logic := '0'; 
signal C_22_S_4_L_7_out : std_logic := '0'; 
signal C_23_S_0_L_0_out : std_logic := '0'; 
signal C_23_S_0_L_1_out : std_logic := '0'; 
signal C_23_S_0_L_2_out : std_logic := '0'; 
signal C_23_S_0_L_3_out : std_logic := '0'; 
signal C_23_S_0_L_4_out : std_logic := '0'; 
signal C_23_S_0_L_5_out : std_logic := '0'; 
signal C_23_S_0_L_6_out : std_logic := '0'; 
signal C_23_S_0_L_7_out : std_logic := '0'; 
signal C_23_S_1_L_0_out : std_logic := '0'; 
signal C_23_S_1_L_1_out : std_logic := '0'; 
signal C_23_S_1_L_2_out : std_logic := '0'; 
signal C_23_S_1_L_3_out : std_logic := '0'; 
signal C_23_S_1_L_4_out : std_logic := '0'; 
signal C_23_S_1_L_5_out : std_logic := '0'; 
signal C_23_S_1_L_6_out : std_logic := '0'; 
signal C_23_S_1_L_7_out : std_logic := '0'; 
signal C_23_S_2_L_0_out : std_logic := '0'; 
signal C_23_S_2_L_1_out : std_logic := '0'; 
signal C_23_S_2_L_2_out : std_logic := '0'; 
signal C_23_S_2_L_3_out : std_logic := '0'; 
signal C_23_S_2_L_4_out : std_logic := '0'; 
signal C_23_S_2_L_5_out : std_logic := '0'; 
signal C_23_S_2_L_6_out : std_logic := '0'; 
signal C_23_S_2_L_7_out : std_logic := '0'; 
signal C_23_S_3_L_0_out : std_logic := '0'; 
signal C_23_S_3_L_1_out : std_logic := '0'; 
signal C_23_S_3_L_2_out : std_logic := '0'; 
signal C_23_S_3_L_3_out : std_logic := '0'; 
signal C_23_S_3_L_4_out : std_logic := '0'; 
signal C_23_S_3_L_5_out : std_logic := '0'; 
signal C_23_S_3_L_6_out : std_logic := '0'; 
signal C_23_S_3_L_7_out : std_logic := '0'; 
signal C_23_S_4_L_0_out : std_logic := '0'; 
signal C_23_S_4_L_1_out : std_logic := '0'; 
signal C_23_S_4_L_2_out : std_logic := '0'; 
signal C_23_S_4_L_3_out : std_logic := '0'; 
signal C_23_S_4_L_4_out : std_logic := '0'; 
signal C_23_S_4_L_5_out : std_logic := '0'; 
signal C_23_S_4_L_6_out : std_logic := '0'; 
signal C_23_S_4_L_7_out : std_logic := '0'; 
signal C_24_S_0_L_0_out : std_logic := '0'; 
signal C_24_S_0_L_1_out : std_logic := '0'; 
signal C_24_S_0_L_2_out : std_logic := '0'; 
signal C_24_S_0_L_3_out : std_logic := '0'; 
signal C_24_S_0_L_4_out : std_logic := '0'; 
signal C_24_S_0_L_5_out : std_logic := '0'; 
signal C_24_S_0_L_6_out : std_logic := '0'; 
signal C_24_S_0_L_7_out : std_logic := '0'; 
signal C_24_S_1_L_0_out : std_logic := '0'; 
signal C_24_S_1_L_1_out : std_logic := '0'; 
signal C_24_S_1_L_2_out : std_logic := '0'; 
signal C_24_S_1_L_3_out : std_logic := '0'; 
signal C_24_S_1_L_4_out : std_logic := '0'; 
signal C_24_S_1_L_5_out : std_logic := '0'; 
signal C_24_S_1_L_6_out : std_logic := '0'; 
signal C_24_S_1_L_7_out : std_logic := '0'; 
signal C_24_S_2_L_0_out : std_logic := '0'; 
signal C_24_S_2_L_1_out : std_logic := '0'; 
signal C_24_S_2_L_2_out : std_logic := '0'; 
signal C_24_S_2_L_3_out : std_logic := '0'; 
signal C_24_S_2_L_4_out : std_logic := '0'; 
signal C_24_S_2_L_5_out : std_logic := '0'; 
signal C_24_S_2_L_6_out : std_logic := '0'; 
signal C_24_S_2_L_7_out : std_logic := '0'; 
signal C_24_S_3_L_0_out : std_logic := '0'; 
signal C_24_S_3_L_1_out : std_logic := '0'; 
signal C_24_S_3_L_2_out : std_logic := '0'; 
signal C_24_S_3_L_3_out : std_logic := '0'; 
signal C_24_S_3_L_4_out : std_logic := '0'; 
signal C_24_S_3_L_5_out : std_logic := '0'; 
signal C_24_S_3_L_6_out : std_logic := '0'; 
signal C_24_S_3_L_7_out : std_logic := '0'; 
signal C_24_S_4_L_0_out : std_logic := '0'; 
signal C_24_S_4_L_1_out : std_logic := '0'; 
signal C_24_S_4_L_2_out : std_logic := '0'; 
signal C_24_S_4_L_3_out : std_logic := '0'; 
signal C_24_S_4_L_4_out : std_logic := '0'; 
signal C_24_S_4_L_5_out : std_logic := '0'; 
signal C_24_S_4_L_6_out : std_logic := '0'; 
signal C_24_S_4_L_7_out : std_logic := '0'; 
signal C_25_S_0_L_0_out : std_logic := '0'; 
signal C_25_S_0_L_1_out : std_logic := '0'; 
signal C_25_S_0_L_2_out : std_logic := '0'; 
signal C_25_S_0_L_3_out : std_logic := '0'; 
signal C_25_S_0_L_4_out : std_logic := '0'; 
signal C_25_S_0_L_5_out : std_logic := '0'; 
signal C_25_S_0_L_6_out : std_logic := '0'; 
signal C_25_S_0_L_7_out : std_logic := '0'; 
signal C_25_S_1_L_0_out : std_logic := '0'; 
signal C_25_S_1_L_1_out : std_logic := '0'; 
signal C_25_S_1_L_2_out : std_logic := '0'; 
signal C_25_S_1_L_3_out : std_logic := '0'; 
signal C_25_S_1_L_4_out : std_logic := '0'; 
signal C_25_S_1_L_5_out : std_logic := '0'; 
signal C_25_S_1_L_6_out : std_logic := '0'; 
signal C_25_S_1_L_7_out : std_logic := '0'; 
signal C_25_S_2_L_0_out : std_logic := '0'; 
signal C_25_S_2_L_1_out : std_logic := '0'; 
signal C_25_S_2_L_2_out : std_logic := '0'; 
signal C_25_S_2_L_3_out : std_logic := '0'; 
signal C_25_S_2_L_4_out : std_logic := '0'; 
signal C_25_S_2_L_5_out : std_logic := '0'; 
signal C_25_S_2_L_6_out : std_logic := '0'; 
signal C_25_S_2_L_7_out : std_logic := '0'; 
signal C_25_S_3_L_0_out : std_logic := '0'; 
signal C_25_S_3_L_1_out : std_logic := '0'; 
signal C_25_S_3_L_2_out : std_logic := '0'; 
signal C_25_S_3_L_3_out : std_logic := '0'; 
signal C_25_S_3_L_4_out : std_logic := '0'; 
signal C_25_S_3_L_5_out : std_logic := '0'; 
signal C_25_S_3_L_6_out : std_logic := '0'; 
signal C_25_S_3_L_7_out : std_logic := '0'; 
signal C_25_S_4_L_0_out : std_logic := '0'; 
signal C_25_S_4_L_1_out : std_logic := '0'; 
signal C_25_S_4_L_2_out : std_logic := '0'; 
signal C_25_S_4_L_3_out : std_logic := '0'; 
signal C_25_S_4_L_4_out : std_logic := '0'; 
signal C_25_S_4_L_5_out : std_logic := '0'; 
signal C_25_S_4_L_6_out : std_logic := '0'; 
signal C_25_S_4_L_7_out : std_logic := '0'; 
signal C_26_S_0_L_0_out : std_logic := '0'; 
signal C_26_S_0_L_1_out : std_logic := '0'; 
signal C_26_S_0_L_2_out : std_logic := '0'; 
signal C_26_S_0_L_3_out : std_logic := '0'; 
signal C_26_S_0_L_4_out : std_logic := '0'; 
signal C_26_S_0_L_5_out : std_logic := '0'; 
signal C_26_S_0_L_6_out : std_logic := '0'; 
signal C_26_S_0_L_7_out : std_logic := '0'; 
signal C_26_S_1_L_0_out : std_logic := '0'; 
signal C_26_S_1_L_1_out : std_logic := '0'; 
signal C_26_S_1_L_2_out : std_logic := '0'; 
signal C_26_S_1_L_3_out : std_logic := '0'; 
signal C_26_S_1_L_4_out : std_logic := '0'; 
signal C_26_S_1_L_5_out : std_logic := '0'; 
signal C_26_S_1_L_6_out : std_logic := '0'; 
signal C_26_S_1_L_7_out : std_logic := '0'; 
signal C_26_S_2_L_0_out : std_logic := '0'; 
signal C_26_S_2_L_1_out : std_logic := '0'; 
signal C_26_S_2_L_2_out : std_logic := '0'; 
signal C_26_S_2_L_3_out : std_logic := '0'; 
signal C_26_S_2_L_4_out : std_logic := '0'; 
signal C_26_S_2_L_5_out : std_logic := '0'; 
signal C_26_S_2_L_6_out : std_logic := '0'; 
signal C_26_S_2_L_7_out : std_logic := '0'; 
signal C_26_S_3_L_0_out : std_logic := '0'; 
signal C_26_S_3_L_1_out : std_logic := '0'; 
signal C_26_S_3_L_2_out : std_logic := '0'; 
signal C_26_S_3_L_3_out : std_logic := '0'; 
signal C_26_S_3_L_4_out : std_logic := '0'; 
signal C_26_S_3_L_5_out : std_logic := '0'; 
signal C_26_S_3_L_6_out : std_logic := '0'; 
signal C_26_S_3_L_7_out : std_logic := '0'; 
signal C_26_S_4_L_0_out : std_logic := '0'; 
signal C_26_S_4_L_1_out : std_logic := '0'; 
signal C_26_S_4_L_2_out : std_logic := '0'; 
signal C_26_S_4_L_3_out : std_logic := '0'; 
signal C_26_S_4_L_4_out : std_logic := '0'; 
signal C_26_S_4_L_5_out : std_logic := '0'; 
signal C_26_S_4_L_6_out : std_logic := '0'; 
signal C_26_S_4_L_7_out : std_logic := '0'; 
signal C_27_S_0_L_0_out : std_logic := '0'; 
signal C_27_S_0_L_1_out : std_logic := '0'; 
signal C_27_S_0_L_2_out : std_logic := '0'; 
signal C_27_S_0_L_3_out : std_logic := '0'; 
signal C_27_S_0_L_4_out : std_logic := '0'; 
signal C_27_S_0_L_5_out : std_logic := '0'; 
signal C_27_S_0_L_6_out : std_logic := '0'; 
signal C_27_S_0_L_7_out : std_logic := '0'; 
signal C_27_S_1_L_0_out : std_logic := '0'; 
signal C_27_S_1_L_1_out : std_logic := '0'; 
signal C_27_S_1_L_2_out : std_logic := '0'; 
signal C_27_S_1_L_3_out : std_logic := '0'; 
signal C_27_S_1_L_4_out : std_logic := '0'; 
signal C_27_S_1_L_5_out : std_logic := '0'; 
signal C_27_S_1_L_6_out : std_logic := '0'; 
signal C_27_S_1_L_7_out : std_logic := '0'; 
signal C_27_S_2_L_0_out : std_logic := '0'; 
signal C_27_S_2_L_1_out : std_logic := '0'; 
signal C_27_S_2_L_2_out : std_logic := '0'; 
signal C_27_S_2_L_3_out : std_logic := '0'; 
signal C_27_S_2_L_4_out : std_logic := '0'; 
signal C_27_S_2_L_5_out : std_logic := '0'; 
signal C_27_S_2_L_6_out : std_logic := '0'; 
signal C_27_S_2_L_7_out : std_logic := '0'; 
signal C_27_S_3_L_0_out : std_logic := '0'; 
signal C_27_S_3_L_1_out : std_logic := '0'; 
signal C_27_S_3_L_2_out : std_logic := '0'; 
signal C_27_S_3_L_3_out : std_logic := '0'; 
signal C_27_S_3_L_4_out : std_logic := '0'; 
signal C_27_S_3_L_5_out : std_logic := '0'; 
signal C_27_S_3_L_6_out : std_logic := '0'; 
signal C_27_S_3_L_7_out : std_logic := '0'; 
signal C_27_S_4_L_0_out : std_logic := '0'; 
signal C_27_S_4_L_1_out : std_logic := '0'; 
signal C_27_S_4_L_2_out : std_logic := '0'; 
signal C_27_S_4_L_3_out : std_logic := '0'; 
signal C_27_S_4_L_4_out : std_logic := '0'; 
signal C_27_S_4_L_5_out : std_logic := '0'; 
signal C_27_S_4_L_6_out : std_logic := '0'; 
signal C_27_S_4_L_7_out : std_logic := '0'; 
signal C_28_S_0_L_0_out : std_logic := '0'; 
signal C_28_S_0_L_1_out : std_logic := '0'; 
signal C_28_S_0_L_2_out : std_logic := '0'; 
signal C_28_S_0_L_3_out : std_logic := '0'; 
signal C_28_S_0_L_4_out : std_logic := '0'; 
signal C_28_S_0_L_5_out : std_logic := '0'; 
signal C_28_S_0_L_6_out : std_logic := '0'; 
signal C_28_S_0_L_7_out : std_logic := '0'; 
signal C_28_S_1_L_0_out : std_logic := '0'; 
signal C_28_S_1_L_1_out : std_logic := '0'; 
signal C_28_S_1_L_2_out : std_logic := '0'; 
signal C_28_S_1_L_3_out : std_logic := '0'; 
signal C_28_S_1_L_4_out : std_logic := '0'; 
signal C_28_S_1_L_5_out : std_logic := '0'; 
signal C_28_S_1_L_6_out : std_logic := '0'; 
signal C_28_S_1_L_7_out : std_logic := '0'; 
signal C_28_S_2_L_0_out : std_logic := '0'; 
signal C_28_S_2_L_1_out : std_logic := '0'; 
signal C_28_S_2_L_2_out : std_logic := '0'; 
signal C_28_S_2_L_3_out : std_logic := '0'; 
signal C_28_S_2_L_4_out : std_logic := '0'; 
signal C_28_S_2_L_5_out : std_logic := '0'; 
signal C_28_S_2_L_6_out : std_logic := '0'; 
signal C_28_S_2_L_7_out : std_logic := '0'; 
signal C_28_S_3_L_0_out : std_logic := '0'; 
signal C_28_S_3_L_1_out : std_logic := '0'; 
signal C_28_S_3_L_2_out : std_logic := '0'; 
signal C_28_S_3_L_3_out : std_logic := '0'; 
signal C_28_S_3_L_4_out : std_logic := '0'; 
signal C_28_S_3_L_5_out : std_logic := '0'; 
signal C_28_S_3_L_6_out : std_logic := '0'; 
signal C_28_S_3_L_7_out : std_logic := '0'; 
signal C_28_S_4_L_0_out : std_logic := '0'; 
signal C_28_S_4_L_1_out : std_logic := '0'; 
signal C_28_S_4_L_2_out : std_logic := '0'; 
signal C_28_S_4_L_3_out : std_logic := '0'; 
signal C_28_S_4_L_4_out : std_logic := '0'; 
signal C_28_S_4_L_5_out : std_logic := '0'; 
signal C_28_S_4_L_6_out : std_logic := '0'; 
signal C_28_S_4_L_7_out : std_logic := '0'; 
signal C_29_S_0_L_0_out : std_logic := '0'; 
signal C_29_S_0_L_1_out : std_logic := '0'; 
signal C_29_S_0_L_2_out : std_logic := '0'; 
signal C_29_S_0_L_3_out : std_logic := '0'; 
signal C_29_S_0_L_4_out : std_logic := '0'; 
signal C_29_S_0_L_5_out : std_logic := '0'; 
signal C_29_S_0_L_6_out : std_logic := '0'; 
signal C_29_S_0_L_7_out : std_logic := '0'; 
signal C_29_S_1_L_0_out : std_logic := '0'; 
signal C_29_S_1_L_1_out : std_logic := '0'; 
signal C_29_S_1_L_2_out : std_logic := '0'; 
signal C_29_S_1_L_3_out : std_logic := '0'; 
signal C_29_S_1_L_4_out : std_logic := '0'; 
signal C_29_S_1_L_5_out : std_logic := '0'; 
signal C_29_S_1_L_6_out : std_logic := '0'; 
signal C_29_S_1_L_7_out : std_logic := '0'; 
signal C_29_S_2_L_0_out : std_logic := '0'; 
signal C_29_S_2_L_1_out : std_logic := '0'; 
signal C_29_S_2_L_2_out : std_logic := '0'; 
signal C_29_S_2_L_3_out : std_logic := '0'; 
signal C_29_S_2_L_4_out : std_logic := '0'; 
signal C_29_S_2_L_5_out : std_logic := '0'; 
signal C_29_S_2_L_6_out : std_logic := '0'; 
signal C_29_S_2_L_7_out : std_logic := '0'; 
signal C_29_S_3_L_0_out : std_logic := '0'; 
signal C_29_S_3_L_1_out : std_logic := '0'; 
signal C_29_S_3_L_2_out : std_logic := '0'; 
signal C_29_S_3_L_3_out : std_logic := '0'; 
signal C_29_S_3_L_4_out : std_logic := '0'; 
signal C_29_S_3_L_5_out : std_logic := '0'; 
signal C_29_S_3_L_6_out : std_logic := '0'; 
signal C_29_S_3_L_7_out : std_logic := '0'; 
signal C_29_S_4_L_0_out : std_logic := '0'; 
signal C_29_S_4_L_1_out : std_logic := '0'; 
signal C_29_S_4_L_2_out : std_logic := '0'; 
signal C_29_S_4_L_3_out : std_logic := '0'; 
signal C_29_S_4_L_4_out : std_logic := '0'; 
signal C_29_S_4_L_5_out : std_logic := '0'; 
signal C_29_S_4_L_6_out : std_logic := '0'; 
signal C_29_S_4_L_7_out : std_logic := '0'; 
signal C_30_S_0_L_0_out : std_logic := '0'; 
signal C_30_S_0_L_1_out : std_logic := '0'; 
signal C_30_S_0_L_2_out : std_logic := '0'; 
signal C_30_S_0_L_3_out : std_logic := '0'; 
signal C_30_S_0_L_4_out : std_logic := '0'; 
signal C_30_S_0_L_5_out : std_logic := '0'; 
signal C_30_S_0_L_6_out : std_logic := '0'; 
signal C_30_S_0_L_7_out : std_logic := '0'; 
signal C_30_S_1_L_0_out : std_logic := '0'; 
signal C_30_S_1_L_1_out : std_logic := '0'; 
signal C_30_S_1_L_2_out : std_logic := '0'; 
signal C_30_S_1_L_3_out : std_logic := '0'; 
signal C_30_S_1_L_4_out : std_logic := '0'; 
signal C_30_S_1_L_5_out : std_logic := '0'; 
signal C_30_S_1_L_6_out : std_logic := '0'; 
signal C_30_S_1_L_7_out : std_logic := '0'; 
signal C_30_S_2_L_0_out : std_logic := '0'; 
signal C_30_S_2_L_1_out : std_logic := '0'; 
signal C_30_S_2_L_2_out : std_logic := '0'; 
signal C_30_S_2_L_3_out : std_logic := '0'; 
signal C_30_S_2_L_4_out : std_logic := '0'; 
signal C_30_S_2_L_5_out : std_logic := '0'; 
signal C_30_S_2_L_6_out : std_logic := '0'; 
signal C_30_S_2_L_7_out : std_logic := '0'; 
signal C_30_S_3_L_0_out : std_logic := '0'; 
signal C_30_S_3_L_1_out : std_logic := '0'; 
signal C_30_S_3_L_2_out : std_logic := '0'; 
signal C_30_S_3_L_3_out : std_logic := '0'; 
signal C_30_S_3_L_4_out : std_logic := '0'; 
signal C_30_S_3_L_5_out : std_logic := '0'; 
signal C_30_S_3_L_6_out : std_logic := '0'; 
signal C_30_S_3_L_7_out : std_logic := '0'; 
signal C_30_S_4_L_0_out : std_logic := '0'; 
signal C_30_S_4_L_1_out : std_logic := '0'; 
signal C_30_S_4_L_2_out : std_logic := '0'; 
signal C_30_S_4_L_3_out : std_logic := '0'; 
signal C_30_S_4_L_4_out : std_logic := '0'; 
signal C_30_S_4_L_5_out : std_logic := '0'; 
signal C_30_S_4_L_6_out : std_logic := '0'; 
signal C_30_S_4_L_7_out : std_logic := '0'; 
signal C_31_S_0_L_0_out : std_logic := '0'; 
signal C_31_S_0_L_1_out : std_logic := '0'; 
signal C_31_S_0_L_2_out : std_logic := '0'; 
signal C_31_S_0_L_3_out : std_logic := '0'; 
signal C_31_S_0_L_4_out : std_logic := '0'; 
signal C_31_S_0_L_5_out : std_logic := '0'; 
signal C_31_S_0_L_6_out : std_logic := '0'; 
signal C_31_S_0_L_7_out : std_logic := '0'; 
signal C_31_S_1_L_0_out : std_logic := '0'; 
signal C_31_S_1_L_1_out : std_logic := '0'; 
signal C_31_S_1_L_2_out : std_logic := '0'; 
signal C_31_S_1_L_3_out : std_logic := '0'; 
signal C_31_S_1_L_4_out : std_logic := '0'; 
signal C_31_S_1_L_5_out : std_logic := '0'; 
signal C_31_S_1_L_6_out : std_logic := '0'; 
signal C_31_S_1_L_7_out : std_logic := '0'; 
signal C_31_S_2_L_0_out : std_logic := '0'; 
signal C_31_S_2_L_1_out : std_logic := '0'; 
signal C_31_S_2_L_2_out : std_logic := '0'; 
signal C_31_S_2_L_3_out : std_logic := '0'; 
signal C_31_S_2_L_4_out : std_logic := '0'; 
signal C_31_S_2_L_5_out : std_logic := '0'; 
signal C_31_S_2_L_6_out : std_logic := '0'; 
signal C_31_S_2_L_7_out : std_logic := '0'; 
signal C_31_S_3_L_0_out : std_logic := '0'; 
signal C_31_S_3_L_1_out : std_logic := '0'; 
signal C_31_S_3_L_2_out : std_logic := '0'; 
signal C_31_S_3_L_3_out : std_logic := '0'; 
signal C_31_S_3_L_4_out : std_logic := '0'; 
signal C_31_S_3_L_5_out : std_logic := '0'; 
signal C_31_S_3_L_6_out : std_logic := '0'; 
signal C_31_S_3_L_7_out : std_logic := '0'; 
signal C_31_S_4_L_0_out : std_logic := '0'; 
signal C_31_S_4_L_1_out : std_logic := '0'; 
signal C_31_S_4_L_2_out : std_logic := '0'; 
signal C_31_S_4_L_3_out : std_logic := '0'; 
signal C_31_S_4_L_4_out : std_logic := '0'; 
signal C_31_S_4_L_5_out : std_logic := '0'; 
signal C_31_S_4_L_6_out : std_logic := '0'; 
signal C_31_S_4_L_7_out : std_logic := '0'; 
signal C_32_S_0_L_0_out : std_logic := '0'; 
signal C_32_S_0_L_1_out : std_logic := '0'; 
signal C_32_S_0_L_2_out : std_logic := '0'; 
signal C_32_S_0_L_3_out : std_logic := '0'; 
signal C_32_S_0_L_4_out : std_logic := '0'; 
signal C_32_S_0_L_5_out : std_logic := '0'; 
signal C_32_S_0_L_6_out : std_logic := '0'; 
signal C_32_S_0_L_7_out : std_logic := '0'; 
signal C_32_S_1_L_0_out : std_logic := '0'; 
signal C_32_S_1_L_1_out : std_logic := '0'; 
signal C_32_S_1_L_2_out : std_logic := '0'; 
signal C_32_S_1_L_3_out : std_logic := '0'; 
signal C_32_S_1_L_4_out : std_logic := '0'; 
signal C_32_S_1_L_5_out : std_logic := '0'; 
signal C_32_S_1_L_6_out : std_logic := '0'; 
signal C_32_S_1_L_7_out : std_logic := '0'; 
signal C_32_S_2_L_0_out : std_logic := '0'; 
signal C_32_S_2_L_1_out : std_logic := '0'; 
signal C_32_S_2_L_2_out : std_logic := '0'; 
signal C_32_S_2_L_3_out : std_logic := '0'; 
signal C_32_S_2_L_4_out : std_logic := '0'; 
signal C_32_S_2_L_5_out : std_logic := '0'; 
signal C_32_S_2_L_6_out : std_logic := '0'; 
signal C_32_S_2_L_7_out : std_logic := '0'; 
signal C_32_S_3_L_0_out : std_logic := '0'; 
signal C_32_S_3_L_1_out : std_logic := '0'; 
signal C_32_S_3_L_2_out : std_logic := '0'; 
signal C_32_S_3_L_3_out : std_logic := '0'; 
signal C_32_S_3_L_4_out : std_logic := '0'; 
signal C_32_S_3_L_5_out : std_logic := '0'; 
signal C_32_S_3_L_6_out : std_logic := '0'; 
signal C_32_S_3_L_7_out : std_logic := '0'; 
signal C_32_S_4_L_0_out : std_logic := '0'; 
signal C_32_S_4_L_1_out : std_logic := '0'; 
signal C_32_S_4_L_2_out : std_logic := '0'; 
signal C_32_S_4_L_3_out : std_logic := '0'; 
signal C_32_S_4_L_4_out : std_logic := '0'; 
signal C_32_S_4_L_5_out : std_logic := '0'; 
signal C_32_S_4_L_6_out : std_logic := '0'; 
signal C_32_S_4_L_7_out : std_logic := '0'; 
signal C_33_S_0_L_0_out : std_logic := '0'; 
signal C_33_S_0_L_1_out : std_logic := '0'; 
signal C_33_S_0_L_2_out : std_logic := '0'; 
signal C_33_S_0_L_3_out : std_logic := '0'; 
signal C_33_S_0_L_4_out : std_logic := '0'; 
signal C_33_S_0_L_5_out : std_logic := '0'; 
signal C_33_S_0_L_6_out : std_logic := '0'; 
signal C_33_S_0_L_7_out : std_logic := '0'; 
signal C_33_S_1_L_0_out : std_logic := '0'; 
signal C_33_S_1_L_1_out : std_logic := '0'; 
signal C_33_S_1_L_2_out : std_logic := '0'; 
signal C_33_S_1_L_3_out : std_logic := '0'; 
signal C_33_S_1_L_4_out : std_logic := '0'; 
signal C_33_S_1_L_5_out : std_logic := '0'; 
signal C_33_S_1_L_6_out : std_logic := '0'; 
signal C_33_S_1_L_7_out : std_logic := '0'; 
signal C_33_S_2_L_0_out : std_logic := '0'; 
signal C_33_S_2_L_1_out : std_logic := '0'; 
signal C_33_S_2_L_2_out : std_logic := '0'; 
signal C_33_S_2_L_3_out : std_logic := '0'; 
signal C_33_S_2_L_4_out : std_logic := '0'; 
signal C_33_S_2_L_5_out : std_logic := '0'; 
signal C_33_S_2_L_6_out : std_logic := '0'; 
signal C_33_S_2_L_7_out : std_logic := '0'; 
signal C_33_S_3_L_0_out : std_logic := '0'; 
signal C_33_S_3_L_1_out : std_logic := '0'; 
signal C_33_S_3_L_2_out : std_logic := '0'; 
signal C_33_S_3_L_3_out : std_logic := '0'; 
signal C_33_S_3_L_4_out : std_logic := '0'; 
signal C_33_S_3_L_5_out : std_logic := '0'; 
signal C_33_S_3_L_6_out : std_logic := '0'; 
signal C_33_S_3_L_7_out : std_logic := '0'; 
signal C_33_S_4_L_0_out : std_logic := '0'; 
signal C_33_S_4_L_1_out : std_logic := '0'; 
signal C_33_S_4_L_2_out : std_logic := '0'; 
signal C_33_S_4_L_3_out : std_logic := '0'; 
signal C_33_S_4_L_4_out : std_logic := '0'; 
signal C_33_S_4_L_5_out : std_logic := '0'; 
signal C_33_S_4_L_6_out : std_logic := '0'; 
signal C_33_S_4_L_7_out : std_logic := '0'; 
signal C_34_S_0_L_0_out : std_logic := '0'; 
signal C_34_S_0_L_1_out : std_logic := '0'; 
signal C_34_S_0_L_2_out : std_logic := '0'; 
signal C_34_S_0_L_3_out : std_logic := '0'; 
signal C_34_S_0_L_4_out : std_logic := '0'; 
signal C_34_S_0_L_5_out : std_logic := '0'; 
signal C_34_S_0_L_6_out : std_logic := '0'; 
signal C_34_S_0_L_7_out : std_logic := '0'; 
signal C_34_S_1_L_0_out : std_logic := '0'; 
signal C_34_S_1_L_1_out : std_logic := '0'; 
signal C_34_S_1_L_2_out : std_logic := '0'; 
signal C_34_S_1_L_3_out : std_logic := '0'; 
signal C_34_S_1_L_4_out : std_logic := '0'; 
signal C_34_S_1_L_5_out : std_logic := '0'; 
signal C_34_S_1_L_6_out : std_logic := '0'; 
signal C_34_S_1_L_7_out : std_logic := '0'; 
signal C_34_S_2_L_0_out : std_logic := '0'; 
signal C_34_S_2_L_1_out : std_logic := '0'; 
signal C_34_S_2_L_2_out : std_logic := '0'; 
signal C_34_S_2_L_3_out : std_logic := '0'; 
signal C_34_S_2_L_4_out : std_logic := '0'; 
signal C_34_S_2_L_5_out : std_logic := '0'; 
signal C_34_S_2_L_6_out : std_logic := '0'; 
signal C_34_S_2_L_7_out : std_logic := '0'; 
signal C_34_S_3_L_0_out : std_logic := '0'; 
signal C_34_S_3_L_1_out : std_logic := '0'; 
signal C_34_S_3_L_2_out : std_logic := '0'; 
signal C_34_S_3_L_3_out : std_logic := '0'; 
signal C_34_S_3_L_4_out : std_logic := '0'; 
signal C_34_S_3_L_5_out : std_logic := '0'; 
signal C_34_S_3_L_6_out : std_logic := '0'; 
signal C_34_S_3_L_7_out : std_logic := '0'; 
signal C_34_S_4_L_0_out : std_logic := '0'; 
signal C_34_S_4_L_1_out : std_logic := '0'; 
signal C_34_S_4_L_2_out : std_logic := '0'; 
signal C_34_S_4_L_3_out : std_logic := '0'; 
signal C_34_S_4_L_4_out : std_logic := '0'; 
signal C_34_S_4_L_5_out : std_logic := '0'; 
signal C_34_S_4_L_6_out : std_logic := '0'; 
signal C_34_S_4_L_7_out : std_logic := '0'; 
signal C_35_S_0_L_0_out : std_logic := '0'; 
signal C_35_S_0_L_1_out : std_logic := '0'; 
signal C_35_S_0_L_2_out : std_logic := '0'; 
signal C_35_S_0_L_3_out : std_logic := '0'; 
signal C_35_S_0_L_4_out : std_logic := '0'; 
signal C_35_S_0_L_5_out : std_logic := '0'; 
signal C_35_S_0_L_6_out : std_logic := '0'; 
signal C_35_S_0_L_7_out : std_logic := '0'; 
signal C_35_S_1_L_0_out : std_logic := '0'; 
signal C_35_S_1_L_1_out : std_logic := '0'; 
signal C_35_S_1_L_2_out : std_logic := '0'; 
signal C_35_S_1_L_3_out : std_logic := '0'; 
signal C_35_S_1_L_4_out : std_logic := '0'; 
signal C_35_S_1_L_5_out : std_logic := '0'; 
signal C_35_S_1_L_6_out : std_logic := '0'; 
signal C_35_S_1_L_7_out : std_logic := '0'; 
signal C_35_S_2_L_0_out : std_logic := '0'; 
signal C_35_S_2_L_1_out : std_logic := '0'; 
signal C_35_S_2_L_2_out : std_logic := '0'; 
signal C_35_S_2_L_3_out : std_logic := '0'; 
signal C_35_S_2_L_4_out : std_logic := '0'; 
signal C_35_S_2_L_5_out : std_logic := '0'; 
signal C_35_S_2_L_6_out : std_logic := '0'; 
signal C_35_S_2_L_7_out : std_logic := '0'; 
signal C_35_S_3_L_0_out : std_logic := '0'; 
signal C_35_S_3_L_1_out : std_logic := '0'; 
signal C_35_S_3_L_2_out : std_logic := '0'; 
signal C_35_S_3_L_3_out : std_logic := '0'; 
signal C_35_S_3_L_4_out : std_logic := '0'; 
signal C_35_S_3_L_5_out : std_logic := '0'; 
signal C_35_S_3_L_6_out : std_logic := '0'; 
signal C_35_S_3_L_7_out : std_logic := '0'; 
signal C_35_S_4_L_0_out : std_logic := '0'; 
signal C_35_S_4_L_1_out : std_logic := '0'; 
signal C_35_S_4_L_2_out : std_logic := '0'; 
signal C_35_S_4_L_3_out : std_logic := '0'; 
signal C_35_S_4_L_4_out : std_logic := '0'; 
signal C_35_S_4_L_5_out : std_logic := '0'; 
signal C_35_S_4_L_6_out : std_logic := '0'; 
signal C_35_S_4_L_7_out : std_logic := '0'; 
signal C_36_S_0_L_0_out : std_logic := '0'; 
signal C_36_S_0_L_1_out : std_logic := '0'; 
signal C_36_S_0_L_2_out : std_logic := '0'; 
signal C_36_S_0_L_3_out : std_logic := '0'; 
signal C_36_S_0_L_4_out : std_logic := '0'; 
signal C_36_S_0_L_5_out : std_logic := '0'; 
signal C_36_S_0_L_6_out : std_logic := '0'; 
signal C_36_S_0_L_7_out : std_logic := '0'; 
signal C_36_S_1_L_0_out : std_logic := '0'; 
signal C_36_S_1_L_1_out : std_logic := '0'; 
signal C_36_S_1_L_2_out : std_logic := '0'; 
signal C_36_S_1_L_3_out : std_logic := '0'; 
signal C_36_S_1_L_4_out : std_logic := '0'; 
signal C_36_S_1_L_5_out : std_logic := '0'; 
signal C_36_S_1_L_6_out : std_logic := '0'; 
signal C_36_S_1_L_7_out : std_logic := '0'; 
signal C_36_S_2_L_0_out : std_logic := '0'; 
signal C_36_S_2_L_1_out : std_logic := '0'; 
signal C_36_S_2_L_2_out : std_logic := '0'; 
signal C_36_S_2_L_3_out : std_logic := '0'; 
signal C_36_S_2_L_4_out : std_logic := '0'; 
signal C_36_S_2_L_5_out : std_logic := '0'; 
signal C_36_S_2_L_6_out : std_logic := '0'; 
signal C_36_S_2_L_7_out : std_logic := '0'; 
signal C_36_S_3_L_0_out : std_logic := '0'; 
signal C_36_S_3_L_1_out : std_logic := '0'; 
signal C_36_S_3_L_2_out : std_logic := '0'; 
signal C_36_S_3_L_3_out : std_logic := '0'; 
signal C_36_S_3_L_4_out : std_logic := '0'; 
signal C_36_S_3_L_5_out : std_logic := '0'; 
signal C_36_S_3_L_6_out : std_logic := '0'; 
signal C_36_S_3_L_7_out : std_logic := '0'; 
signal C_36_S_4_L_0_out : std_logic := '0'; 
signal C_36_S_4_L_1_out : std_logic := '0'; 
signal C_36_S_4_L_2_out : std_logic := '0'; 
signal C_36_S_4_L_3_out : std_logic := '0'; 
signal C_36_S_4_L_4_out : std_logic := '0'; 
signal C_36_S_4_L_5_out : std_logic := '0'; 
signal C_36_S_4_L_6_out : std_logic := '0'; 
signal C_36_S_4_L_7_out : std_logic := '0'; 
signal C_37_S_0_L_0_out : std_logic := '0'; 
signal C_37_S_0_L_1_out : std_logic := '0'; 
signal C_37_S_0_L_2_out : std_logic := '0'; 
signal C_37_S_0_L_3_out : std_logic := '0'; 
signal C_37_S_0_L_4_out : std_logic := '0'; 
signal C_37_S_0_L_5_out : std_logic := '0'; 
signal C_37_S_0_L_6_out : std_logic := '0'; 
signal C_37_S_0_L_7_out : std_logic := '0'; 
signal C_37_S_1_L_0_out : std_logic := '0'; 
signal C_37_S_1_L_1_out : std_logic := '0'; 
signal C_37_S_1_L_2_out : std_logic := '0'; 
signal C_37_S_1_L_3_out : std_logic := '0'; 
signal C_37_S_1_L_4_out : std_logic := '0'; 
signal C_37_S_1_L_5_out : std_logic := '0'; 
signal C_37_S_1_L_6_out : std_logic := '0'; 
signal C_37_S_1_L_7_out : std_logic := '0'; 
signal C_37_S_2_L_0_out : std_logic := '0'; 
signal C_37_S_2_L_1_out : std_logic := '0'; 
signal C_37_S_2_L_2_out : std_logic := '0'; 
signal C_37_S_2_L_3_out : std_logic := '0'; 
signal C_37_S_2_L_4_out : std_logic := '0'; 
signal C_37_S_2_L_5_out : std_logic := '0'; 
signal C_37_S_2_L_6_out : std_logic := '0'; 
signal C_37_S_2_L_7_out : std_logic := '0'; 
signal C_37_S_3_L_0_out : std_logic := '0'; 
signal C_37_S_3_L_1_out : std_logic := '0'; 
signal C_37_S_3_L_2_out : std_logic := '0'; 
signal C_37_S_3_L_3_out : std_logic := '0'; 
signal C_37_S_3_L_4_out : std_logic := '0'; 
signal C_37_S_3_L_5_out : std_logic := '0'; 
signal C_37_S_3_L_6_out : std_logic := '0'; 
signal C_37_S_3_L_7_out : std_logic := '0'; 
signal C_37_S_4_L_0_out : std_logic := '0'; 
signal C_37_S_4_L_1_out : std_logic := '0'; 
signal C_37_S_4_L_2_out : std_logic := '0'; 
signal C_37_S_4_L_3_out : std_logic := '0'; 
signal C_37_S_4_L_4_out : std_logic := '0'; 
signal C_37_S_4_L_5_out : std_logic := '0'; 
signal C_37_S_4_L_6_out : std_logic := '0'; 
signal C_37_S_4_L_7_out : std_logic := '0'; 
signal C_38_S_0_L_0_out : std_logic := '0'; 
signal C_38_S_0_L_1_out : std_logic := '0'; 
signal C_38_S_0_L_2_out : std_logic := '0'; 
signal C_38_S_0_L_3_out : std_logic := '0'; 
signal C_38_S_0_L_4_out : std_logic := '0'; 
signal C_38_S_0_L_5_out : std_logic := '0'; 
signal C_38_S_0_L_6_out : std_logic := '0'; 
signal C_38_S_0_L_7_out : std_logic := '0'; 
signal C_38_S_1_L_0_out : std_logic := '0'; 
signal C_38_S_1_L_1_out : std_logic := '0'; 
signal C_38_S_1_L_2_out : std_logic := '0'; 
signal C_38_S_1_L_3_out : std_logic := '0'; 
signal C_38_S_1_L_4_out : std_logic := '0'; 
signal C_38_S_1_L_5_out : std_logic := '0'; 
signal C_38_S_1_L_6_out : std_logic := '0'; 
signal C_38_S_1_L_7_out : std_logic := '0'; 
signal C_38_S_2_L_0_out : std_logic := '0'; 
signal C_38_S_2_L_1_out : std_logic := '0'; 
signal C_38_S_2_L_2_out : std_logic := '0'; 
signal C_38_S_2_L_3_out : std_logic := '0'; 
signal C_38_S_2_L_4_out : std_logic := '0'; 
signal C_38_S_2_L_5_out : std_logic := '0'; 
signal C_38_S_2_L_6_out : std_logic := '0'; 
signal C_38_S_2_L_7_out : std_logic := '0'; 
signal C_38_S_3_L_0_out : std_logic := '0'; 
signal C_38_S_3_L_1_out : std_logic := '0'; 
signal C_38_S_3_L_2_out : std_logic := '0'; 
signal C_38_S_3_L_3_out : std_logic := '0'; 
signal C_38_S_3_L_4_out : std_logic := '0'; 
signal C_38_S_3_L_5_out : std_logic := '0'; 
signal C_38_S_3_L_6_out : std_logic := '0'; 
signal C_38_S_3_L_7_out : std_logic := '0'; 
signal C_38_S_4_L_0_out : std_logic := '0'; 
signal C_38_S_4_L_1_out : std_logic := '0'; 
signal C_38_S_4_L_2_out : std_logic := '0'; 
signal C_38_S_4_L_3_out : std_logic := '0'; 
signal C_38_S_4_L_4_out : std_logic := '0'; 
signal C_38_S_4_L_5_out : std_logic := '0'; 
signal C_38_S_4_L_6_out : std_logic := '0'; 
signal C_38_S_4_L_7_out : std_logic := '0'; 
signal C_39_S_0_L_0_out : std_logic := '0'; 
signal C_39_S_0_L_1_out : std_logic := '0'; 
signal C_39_S_0_L_2_out : std_logic := '0'; 
signal C_39_S_0_L_3_out : std_logic := '0'; 
signal C_39_S_0_L_4_out : std_logic := '0'; 
signal C_39_S_0_L_5_out : std_logic := '0'; 
signal C_39_S_0_L_6_out : std_logic := '0'; 
signal C_39_S_0_L_7_out : std_logic := '0'; 
signal C_39_S_1_L_0_out : std_logic := '0'; 
signal C_39_S_1_L_1_out : std_logic := '0'; 
signal C_39_S_1_L_2_out : std_logic := '0'; 
signal C_39_S_1_L_3_out : std_logic := '0'; 
signal C_39_S_1_L_4_out : std_logic := '0'; 
signal C_39_S_1_L_5_out : std_logic := '0'; 
signal C_39_S_1_L_6_out : std_logic := '0'; 
signal C_39_S_1_L_7_out : std_logic := '0'; 
signal C_39_S_2_L_0_out : std_logic := '0'; 
signal C_39_S_2_L_1_out : std_logic := '0'; 
signal C_39_S_2_L_2_out : std_logic := '0'; 
signal C_39_S_2_L_3_out : std_logic := '0'; 
signal C_39_S_2_L_4_out : std_logic := '0'; 
signal C_39_S_2_L_5_out : std_logic := '0'; 
signal C_39_S_2_L_6_out : std_logic := '0'; 
signal C_39_S_2_L_7_out : std_logic := '0'; 
signal C_39_S_3_L_0_out : std_logic := '0'; 
signal C_39_S_3_L_1_out : std_logic := '0'; 
signal C_39_S_3_L_2_out : std_logic := '0'; 
signal C_39_S_3_L_3_out : std_logic := '0'; 
signal C_39_S_3_L_4_out : std_logic := '0'; 
signal C_39_S_3_L_5_out : std_logic := '0'; 
signal C_39_S_3_L_6_out : std_logic := '0'; 
signal C_39_S_3_L_7_out : std_logic := '0'; 
signal C_39_S_4_L_0_out : std_logic := '0'; 
signal C_39_S_4_L_1_out : std_logic := '0'; 
signal C_39_S_4_L_2_out : std_logic := '0'; 
signal C_39_S_4_L_3_out : std_logic := '0'; 
signal C_39_S_4_L_4_out : std_logic := '0'; 
signal C_39_S_4_L_5_out : std_logic := '0'; 
signal C_39_S_4_L_6_out : std_logic := '0'; 
signal C_39_S_4_L_7_out : std_logic := '0'; 
signal C_40_S_0_L_0_out : std_logic := '0'; 
signal C_40_S_0_L_1_out : std_logic := '0'; 
signal C_40_S_0_L_2_out : std_logic := '0'; 
signal C_40_S_0_L_3_out : std_logic := '0'; 
signal C_40_S_0_L_4_out : std_logic := '0'; 
signal C_40_S_0_L_5_out : std_logic := '0'; 
signal C_40_S_0_L_6_out : std_logic := '0'; 
signal C_40_S_0_L_7_out : std_logic := '0'; 
signal C_40_S_1_L_0_out : std_logic := '0'; 
signal C_40_S_1_L_1_out : std_logic := '0'; 
signal C_40_S_1_L_2_out : std_logic := '0'; 
signal C_40_S_1_L_3_out : std_logic := '0'; 
signal C_40_S_1_L_4_out : std_logic := '0'; 
signal C_40_S_1_L_5_out : std_logic := '0'; 
signal C_40_S_1_L_6_out : std_logic := '0'; 
signal C_40_S_1_L_7_out : std_logic := '0'; 
signal C_40_S_2_L_0_out : std_logic := '0'; 
signal C_40_S_2_L_1_out : std_logic := '0'; 
signal C_40_S_2_L_2_out : std_logic := '0'; 
signal C_40_S_2_L_3_out : std_logic := '0'; 
signal C_40_S_2_L_4_out : std_logic := '0'; 
signal C_40_S_2_L_5_out : std_logic := '0'; 
signal C_40_S_2_L_6_out : std_logic := '0'; 
signal C_40_S_2_L_7_out : std_logic := '0'; 
signal C_40_S_3_L_0_out : std_logic := '0'; 
signal C_40_S_3_L_1_out : std_logic := '0'; 
signal C_40_S_3_L_2_out : std_logic := '0'; 
signal C_40_S_3_L_3_out : std_logic := '0'; 
signal C_40_S_3_L_4_out : std_logic := '0'; 
signal C_40_S_3_L_5_out : std_logic := '0'; 
signal C_40_S_3_L_6_out : std_logic := '0'; 
signal C_40_S_3_L_7_out : std_logic := '0'; 
signal C_40_S_4_L_0_out : std_logic := '0'; 
signal C_40_S_4_L_1_out : std_logic := '0'; 
signal C_40_S_4_L_2_out : std_logic := '0'; 
signal C_40_S_4_L_3_out : std_logic := '0'; 
signal C_40_S_4_L_4_out : std_logic := '0'; 
signal C_40_S_4_L_5_out : std_logic := '0'; 
signal C_40_S_4_L_6_out : std_logic := '0'; 
signal C_40_S_4_L_7_out : std_logic := '0'; 
signal C_41_S_0_L_0_out : std_logic := '0'; 
signal C_41_S_0_L_1_out : std_logic := '0'; 
signal C_41_S_0_L_2_out : std_logic := '0'; 
signal C_41_S_0_L_3_out : std_logic := '0'; 
signal C_41_S_0_L_4_out : std_logic := '0'; 
signal C_41_S_0_L_5_out : std_logic := '0'; 
signal C_41_S_0_L_6_out : std_logic := '0'; 
signal C_41_S_0_L_7_out : std_logic := '0'; 
signal C_41_S_1_L_0_out : std_logic := '0'; 
signal C_41_S_1_L_1_out : std_logic := '0'; 
signal C_41_S_1_L_2_out : std_logic := '0'; 
signal C_41_S_1_L_3_out : std_logic := '0'; 
signal C_41_S_1_L_4_out : std_logic := '0'; 
signal C_41_S_1_L_5_out : std_logic := '0'; 
signal C_41_S_1_L_6_out : std_logic := '0'; 
signal C_41_S_1_L_7_out : std_logic := '0'; 
signal C_41_S_2_L_0_out : std_logic := '0'; 
signal C_41_S_2_L_1_out : std_logic := '0'; 
signal C_41_S_2_L_2_out : std_logic := '0'; 
signal C_41_S_2_L_3_out : std_logic := '0'; 
signal C_41_S_2_L_4_out : std_logic := '0'; 
signal C_41_S_2_L_5_out : std_logic := '0'; 
signal C_41_S_2_L_6_out : std_logic := '0'; 
signal C_41_S_2_L_7_out : std_logic := '0'; 
signal C_41_S_3_L_0_out : std_logic := '0'; 
signal C_41_S_3_L_1_out : std_logic := '0'; 
signal C_41_S_3_L_2_out : std_logic := '0'; 
signal C_41_S_3_L_3_out : std_logic := '0'; 
signal C_41_S_3_L_4_out : std_logic := '0'; 
signal C_41_S_3_L_5_out : std_logic := '0'; 
signal C_41_S_3_L_6_out : std_logic := '0'; 
signal C_41_S_3_L_7_out : std_logic := '0'; 
signal C_41_S_4_L_0_out : std_logic := '0'; 
signal C_41_S_4_L_1_out : std_logic := '0'; 
signal C_41_S_4_L_2_out : std_logic := '0'; 
signal C_41_S_4_L_3_out : std_logic := '0'; 
signal C_41_S_4_L_4_out : std_logic := '0'; 
signal C_41_S_4_L_5_out : std_logic := '0'; 
signal C_41_S_4_L_6_out : std_logic := '0'; 
signal C_41_S_4_L_7_out : std_logic := '0'; 
signal C_42_S_0_L_0_out : std_logic := '0'; 
signal C_42_S_0_L_1_out : std_logic := '0'; 
signal C_42_S_0_L_2_out : std_logic := '0'; 
signal C_42_S_0_L_3_out : std_logic := '0'; 
signal C_42_S_0_L_4_out : std_logic := '0'; 
signal C_42_S_0_L_5_out : std_logic := '0'; 
signal C_42_S_0_L_6_out : std_logic := '0'; 
signal C_42_S_0_L_7_out : std_logic := '0'; 
signal C_42_S_1_L_0_out : std_logic := '0'; 
signal C_42_S_1_L_1_out : std_logic := '0'; 
signal C_42_S_1_L_2_out : std_logic := '0'; 
signal C_42_S_1_L_3_out : std_logic := '0'; 
signal C_42_S_1_L_4_out : std_logic := '0'; 
signal C_42_S_1_L_5_out : std_logic := '0'; 
signal C_42_S_1_L_6_out : std_logic := '0'; 
signal C_42_S_1_L_7_out : std_logic := '0'; 
signal C_42_S_2_L_0_out : std_logic := '0'; 
signal C_42_S_2_L_1_out : std_logic := '0'; 
signal C_42_S_2_L_2_out : std_logic := '0'; 
signal C_42_S_2_L_3_out : std_logic := '0'; 
signal C_42_S_2_L_4_out : std_logic := '0'; 
signal C_42_S_2_L_5_out : std_logic := '0'; 
signal C_42_S_2_L_6_out : std_logic := '0'; 
signal C_42_S_2_L_7_out : std_logic := '0'; 
signal C_42_S_3_L_0_out : std_logic := '0'; 
signal C_42_S_3_L_1_out : std_logic := '0'; 
signal C_42_S_3_L_2_out : std_logic := '0'; 
signal C_42_S_3_L_3_out : std_logic := '0'; 
signal C_42_S_3_L_4_out : std_logic := '0'; 
signal C_42_S_3_L_5_out : std_logic := '0'; 
signal C_42_S_3_L_6_out : std_logic := '0'; 
signal C_42_S_3_L_7_out : std_logic := '0'; 
signal C_42_S_4_L_0_out : std_logic := '0'; 
signal C_42_S_4_L_1_out : std_logic := '0'; 
signal C_42_S_4_L_2_out : std_logic := '0'; 
signal C_42_S_4_L_3_out : std_logic := '0'; 
signal C_42_S_4_L_4_out : std_logic := '0'; 
signal C_42_S_4_L_5_out : std_logic := '0'; 
signal C_42_S_4_L_6_out : std_logic := '0'; 
signal C_42_S_4_L_7_out : std_logic := '0'; 
signal C_43_S_0_L_0_out : std_logic := '0'; 
signal C_43_S_0_L_1_out : std_logic := '0'; 
signal C_43_S_0_L_2_out : std_logic := '0'; 
signal C_43_S_0_L_3_out : std_logic := '0'; 
signal C_43_S_0_L_4_out : std_logic := '0'; 
signal C_43_S_0_L_5_out : std_logic := '0'; 
signal C_43_S_0_L_6_out : std_logic := '0'; 
signal C_43_S_0_L_7_out : std_logic := '0'; 
signal C_43_S_1_L_0_out : std_logic := '0'; 
signal C_43_S_1_L_1_out : std_logic := '0'; 
signal C_43_S_1_L_2_out : std_logic := '0'; 
signal C_43_S_1_L_3_out : std_logic := '0'; 
signal C_43_S_1_L_4_out : std_logic := '0'; 
signal C_43_S_1_L_5_out : std_logic := '0'; 
signal C_43_S_1_L_6_out : std_logic := '0'; 
signal C_43_S_1_L_7_out : std_logic := '0'; 
signal C_43_S_2_L_0_out : std_logic := '0'; 
signal C_43_S_2_L_1_out : std_logic := '0'; 
signal C_43_S_2_L_2_out : std_logic := '0'; 
signal C_43_S_2_L_3_out : std_logic := '0'; 
signal C_43_S_2_L_4_out : std_logic := '0'; 
signal C_43_S_2_L_5_out : std_logic := '0'; 
signal C_43_S_2_L_6_out : std_logic := '0'; 
signal C_43_S_2_L_7_out : std_logic := '0'; 
signal C_43_S_3_L_0_out : std_logic := '0'; 
signal C_43_S_3_L_1_out : std_logic := '0'; 
signal C_43_S_3_L_2_out : std_logic := '0'; 
signal C_43_S_3_L_3_out : std_logic := '0'; 
signal C_43_S_3_L_4_out : std_logic := '0'; 
signal C_43_S_3_L_5_out : std_logic := '0'; 
signal C_43_S_3_L_6_out : std_logic := '0'; 
signal C_43_S_3_L_7_out : std_logic := '0'; 
signal C_43_S_4_L_0_out : std_logic := '0'; 
signal C_43_S_4_L_1_out : std_logic := '0'; 
signal C_43_S_4_L_2_out : std_logic := '0'; 
signal C_43_S_4_L_3_out : std_logic := '0'; 
signal C_43_S_4_L_4_out : std_logic := '0'; 
signal C_43_S_4_L_5_out : std_logic := '0'; 
signal C_43_S_4_L_6_out : std_logic := '0'; 
signal C_43_S_4_L_7_out : std_logic := '0'; 
signal C_44_S_0_L_0_out : std_logic := '0'; 
signal C_44_S_0_L_1_out : std_logic := '0'; 
signal C_44_S_0_L_2_out : std_logic := '0'; 
signal C_44_S_0_L_3_out : std_logic := '0'; 
signal C_44_S_0_L_4_out : std_logic := '0'; 
signal C_44_S_0_L_5_out : std_logic := '0'; 
signal C_44_S_0_L_6_out : std_logic := '0'; 
signal C_44_S_0_L_7_out : std_logic := '0'; 
signal C_44_S_1_L_0_out : std_logic := '0'; 
signal C_44_S_1_L_1_out : std_logic := '0'; 
signal C_44_S_1_L_2_out : std_logic := '0'; 
signal C_44_S_1_L_3_out : std_logic := '0'; 
signal C_44_S_1_L_4_out : std_logic := '0'; 
signal C_44_S_1_L_5_out : std_logic := '0'; 
signal C_44_S_1_L_6_out : std_logic := '0'; 
signal C_44_S_1_L_7_out : std_logic := '0'; 
signal C_44_S_2_L_0_out : std_logic := '0'; 
signal C_44_S_2_L_1_out : std_logic := '0'; 
signal C_44_S_2_L_2_out : std_logic := '0'; 
signal C_44_S_2_L_3_out : std_logic := '0'; 
signal C_44_S_2_L_4_out : std_logic := '0'; 
signal C_44_S_2_L_5_out : std_logic := '0'; 
signal C_44_S_2_L_6_out : std_logic := '0'; 
signal C_44_S_2_L_7_out : std_logic := '0'; 
signal C_44_S_3_L_0_out : std_logic := '0'; 
signal C_44_S_3_L_1_out : std_logic := '0'; 
signal C_44_S_3_L_2_out : std_logic := '0'; 
signal C_44_S_3_L_3_out : std_logic := '0'; 
signal C_44_S_3_L_4_out : std_logic := '0'; 
signal C_44_S_3_L_5_out : std_logic := '0'; 
signal C_44_S_3_L_6_out : std_logic := '0'; 
signal C_44_S_3_L_7_out : std_logic := '0'; 
signal C_44_S_4_L_0_out : std_logic := '0'; 
signal C_44_S_4_L_1_out : std_logic := '0'; 
signal C_44_S_4_L_2_out : std_logic := '0'; 
signal C_44_S_4_L_3_out : std_logic := '0'; 
signal C_44_S_4_L_4_out : std_logic := '0'; 
signal C_44_S_4_L_5_out : std_logic := '0'; 
signal C_44_S_4_L_6_out : std_logic := '0'; 
signal C_44_S_4_L_7_out : std_logic := '0'; 
signal C_45_S_0_L_0_out : std_logic := '0'; 
signal C_45_S_0_L_1_out : std_logic := '0'; 
signal C_45_S_0_L_2_out : std_logic := '0'; 
signal C_45_S_0_L_3_out : std_logic := '0'; 
signal C_45_S_0_L_4_out : std_logic := '0'; 
signal C_45_S_0_L_5_out : std_logic := '0'; 
signal C_45_S_0_L_6_out : std_logic := '0'; 
signal C_45_S_0_L_7_out : std_logic := '0'; 
signal C_45_S_1_L_0_out : std_logic := '0'; 
signal C_45_S_1_L_1_out : std_logic := '0'; 
signal C_45_S_1_L_2_out : std_logic := '0'; 
signal C_45_S_1_L_3_out : std_logic := '0'; 
signal C_45_S_1_L_4_out : std_logic := '0'; 
signal C_45_S_1_L_5_out : std_logic := '0'; 
signal C_45_S_1_L_6_out : std_logic := '0'; 
signal C_45_S_1_L_7_out : std_logic := '0'; 
signal C_45_S_2_L_0_out : std_logic := '0'; 
signal C_45_S_2_L_1_out : std_logic := '0'; 
signal C_45_S_2_L_2_out : std_logic := '0'; 
signal C_45_S_2_L_3_out : std_logic := '0'; 
signal C_45_S_2_L_4_out : std_logic := '0'; 
signal C_45_S_2_L_5_out : std_logic := '0'; 
signal C_45_S_2_L_6_out : std_logic := '0'; 
signal C_45_S_2_L_7_out : std_logic := '0'; 
signal C_45_S_3_L_0_out : std_logic := '0'; 
signal C_45_S_3_L_1_out : std_logic := '0'; 
signal C_45_S_3_L_2_out : std_logic := '0'; 
signal C_45_S_3_L_3_out : std_logic := '0'; 
signal C_45_S_3_L_4_out : std_logic := '0'; 
signal C_45_S_3_L_5_out : std_logic := '0'; 
signal C_45_S_3_L_6_out : std_logic := '0'; 
signal C_45_S_3_L_7_out : std_logic := '0'; 
signal C_45_S_4_L_0_out : std_logic := '0'; 
signal C_45_S_4_L_1_out : std_logic := '0'; 
signal C_45_S_4_L_2_out : std_logic := '0'; 
signal C_45_S_4_L_3_out : std_logic := '0'; 
signal C_45_S_4_L_4_out : std_logic := '0'; 
signal C_45_S_4_L_5_out : std_logic := '0'; 
signal C_45_S_4_L_6_out : std_logic := '0'; 
signal C_45_S_4_L_7_out : std_logic := '0'; 
signal C_46_S_0_L_0_out : std_logic := '0'; 
signal C_46_S_0_L_1_out : std_logic := '0'; 
signal C_46_S_0_L_2_out : std_logic := '0'; 
signal C_46_S_0_L_3_out : std_logic := '0'; 
signal C_46_S_0_L_4_out : std_logic := '0'; 
signal C_46_S_0_L_5_out : std_logic := '0'; 
signal C_46_S_0_L_6_out : std_logic := '0'; 
signal C_46_S_0_L_7_out : std_logic := '0'; 
signal C_46_S_1_L_0_out : std_logic := '0'; 
signal C_46_S_1_L_1_out : std_logic := '0'; 
signal C_46_S_1_L_2_out : std_logic := '0'; 
signal C_46_S_1_L_3_out : std_logic := '0'; 
signal C_46_S_1_L_4_out : std_logic := '0'; 
signal C_46_S_1_L_5_out : std_logic := '0'; 
signal C_46_S_1_L_6_out : std_logic := '0'; 
signal C_46_S_1_L_7_out : std_logic := '0'; 
signal C_46_S_2_L_0_out : std_logic := '0'; 
signal C_46_S_2_L_1_out : std_logic := '0'; 
signal C_46_S_2_L_2_out : std_logic := '0'; 
signal C_46_S_2_L_3_out : std_logic := '0'; 
signal C_46_S_2_L_4_out : std_logic := '0'; 
signal C_46_S_2_L_5_out : std_logic := '0'; 
signal C_46_S_2_L_6_out : std_logic := '0'; 
signal C_46_S_2_L_7_out : std_logic := '0'; 
signal C_46_S_3_L_0_out : std_logic := '0'; 
signal C_46_S_3_L_1_out : std_logic := '0'; 
signal C_46_S_3_L_2_out : std_logic := '0'; 
signal C_46_S_3_L_3_out : std_logic := '0'; 
signal C_46_S_3_L_4_out : std_logic := '0'; 
signal C_46_S_3_L_5_out : std_logic := '0'; 
signal C_46_S_3_L_6_out : std_logic := '0'; 
signal C_46_S_3_L_7_out : std_logic := '0'; 
signal C_46_S_4_L_0_out : std_logic := '0'; 
signal C_46_S_4_L_1_out : std_logic := '0'; 
signal C_46_S_4_L_2_out : std_logic := '0'; 
signal C_46_S_4_L_3_out : std_logic := '0'; 
signal C_46_S_4_L_4_out : std_logic := '0'; 
signal C_46_S_4_L_5_out : std_logic := '0'; 
signal C_46_S_4_L_6_out : std_logic := '0'; 
signal C_46_S_4_L_7_out : std_logic := '0'; 
signal C_47_S_0_L_0_out : std_logic := '0'; 
signal C_47_S_0_L_1_out : std_logic := '0'; 
signal C_47_S_0_L_2_out : std_logic := '0'; 
signal C_47_S_0_L_3_out : std_logic := '0'; 
signal C_47_S_0_L_4_out : std_logic := '0'; 
signal C_47_S_0_L_5_out : std_logic := '0'; 
signal C_47_S_0_L_6_out : std_logic := '0'; 
signal C_47_S_0_L_7_out : std_logic := '0'; 
signal C_47_S_1_L_0_out : std_logic := '0'; 
signal C_47_S_1_L_1_out : std_logic := '0'; 
signal C_47_S_1_L_2_out : std_logic := '0'; 
signal C_47_S_1_L_3_out : std_logic := '0'; 
signal C_47_S_1_L_4_out : std_logic := '0'; 
signal C_47_S_1_L_5_out : std_logic := '0'; 
signal C_47_S_1_L_6_out : std_logic := '0'; 
signal C_47_S_1_L_7_out : std_logic := '0'; 
signal C_47_S_2_L_0_out : std_logic := '0'; 
signal C_47_S_2_L_1_out : std_logic := '0'; 
signal C_47_S_2_L_2_out : std_logic := '0'; 
signal C_47_S_2_L_3_out : std_logic := '0'; 
signal C_47_S_2_L_4_out : std_logic := '0'; 
signal C_47_S_2_L_5_out : std_logic := '0'; 
signal C_47_S_2_L_6_out : std_logic := '0'; 
signal C_47_S_2_L_7_out : std_logic := '0'; 
signal C_47_S_3_L_0_out : std_logic := '0'; 
signal C_47_S_3_L_1_out : std_logic := '0'; 
signal C_47_S_3_L_2_out : std_logic := '0'; 
signal C_47_S_3_L_3_out : std_logic := '0'; 
signal C_47_S_3_L_4_out : std_logic := '0'; 
signal C_47_S_3_L_5_out : std_logic := '0'; 
signal C_47_S_3_L_6_out : std_logic := '0'; 
signal C_47_S_3_L_7_out : std_logic := '0'; 
signal C_47_S_4_L_0_out : std_logic := '0'; 
signal C_47_S_4_L_1_out : std_logic := '0'; 
signal C_47_S_4_L_2_out : std_logic := '0'; 
signal C_47_S_4_L_3_out : std_logic := '0'; 
signal C_47_S_4_L_4_out : std_logic := '0'; 
signal C_47_S_4_L_5_out : std_logic := '0'; 
signal C_47_S_4_L_6_out : std_logic := '0'; 
signal C_47_S_4_L_7_out : std_logic := '0'; 
signal C_48_S_0_L_0_out : std_logic := '0'; 
signal C_48_S_0_L_1_out : std_logic := '0'; 
signal C_48_S_0_L_2_out : std_logic := '0'; 
signal C_48_S_0_L_3_out : std_logic := '0'; 
signal C_48_S_0_L_4_out : std_logic := '0'; 
signal C_48_S_0_L_5_out : std_logic := '0'; 
signal C_48_S_0_L_6_out : std_logic := '0'; 
signal C_48_S_0_L_7_out : std_logic := '0'; 
signal C_48_S_1_L_0_out : std_logic := '0'; 
signal C_48_S_1_L_1_out : std_logic := '0'; 
signal C_48_S_1_L_2_out : std_logic := '0'; 
signal C_48_S_1_L_3_out : std_logic := '0'; 
signal C_48_S_1_L_4_out : std_logic := '0'; 
signal C_48_S_1_L_5_out : std_logic := '0'; 
signal C_48_S_1_L_6_out : std_logic := '0'; 
signal C_48_S_1_L_7_out : std_logic := '0'; 
signal C_48_S_2_L_0_out : std_logic := '0'; 
signal C_48_S_2_L_1_out : std_logic := '0'; 
signal C_48_S_2_L_2_out : std_logic := '0'; 
signal C_48_S_2_L_3_out : std_logic := '0'; 
signal C_48_S_2_L_4_out : std_logic := '0'; 
signal C_48_S_2_L_5_out : std_logic := '0'; 
signal C_48_S_2_L_6_out : std_logic := '0'; 
signal C_48_S_2_L_7_out : std_logic := '0'; 
signal C_48_S_3_L_0_out : std_logic := '0'; 
signal C_48_S_3_L_1_out : std_logic := '0'; 
signal C_48_S_3_L_2_out : std_logic := '0'; 
signal C_48_S_3_L_3_out : std_logic := '0'; 
signal C_48_S_3_L_4_out : std_logic := '0'; 
signal C_48_S_3_L_5_out : std_logic := '0'; 
signal C_48_S_3_L_6_out : std_logic := '0'; 
signal C_48_S_3_L_7_out : std_logic := '0'; 
signal C_48_S_4_L_0_out : std_logic := '0'; 
signal C_48_S_4_L_1_out : std_logic := '0'; 
signal C_48_S_4_L_2_out : std_logic := '0'; 
signal C_48_S_4_L_3_out : std_logic := '0'; 
signal C_48_S_4_L_4_out : std_logic := '0'; 
signal C_48_S_4_L_5_out : std_logic := '0'; 
signal C_48_S_4_L_6_out : std_logic := '0'; 
signal C_48_S_4_L_7_out : std_logic := '0'; 
signal C_49_S_0_L_0_out : std_logic := '0'; 
signal C_49_S_0_L_1_out : std_logic := '0'; 
signal C_49_S_0_L_2_out : std_logic := '0'; 
signal C_49_S_0_L_3_out : std_logic := '0'; 
signal C_49_S_0_L_4_out : std_logic := '0'; 
signal C_49_S_0_L_5_out : std_logic := '0'; 
signal C_49_S_0_L_6_out : std_logic := '0'; 
signal C_49_S_0_L_7_out : std_logic := '0'; 
signal C_49_S_1_L_0_out : std_logic := '0'; 
signal C_49_S_1_L_1_out : std_logic := '0'; 
signal C_49_S_1_L_2_out : std_logic := '0'; 
signal C_49_S_1_L_3_out : std_logic := '0'; 
signal C_49_S_1_L_4_out : std_logic := '0'; 
signal C_49_S_1_L_5_out : std_logic := '0'; 
signal C_49_S_1_L_6_out : std_logic := '0'; 
signal C_49_S_1_L_7_out : std_logic := '0'; 
signal C_49_S_2_L_0_out : std_logic := '0'; 
signal C_49_S_2_L_1_out : std_logic := '0'; 
signal C_49_S_2_L_2_out : std_logic := '0'; 
signal C_49_S_2_L_3_out : std_logic := '0'; 
signal C_49_S_2_L_4_out : std_logic := '0'; 
signal C_49_S_2_L_5_out : std_logic := '0'; 
signal C_49_S_2_L_6_out : std_logic := '0'; 
signal C_49_S_2_L_7_out : std_logic := '0'; 
signal C_49_S_3_L_0_out : std_logic := '0'; 
signal C_49_S_3_L_1_out : std_logic := '0'; 
signal C_49_S_3_L_2_out : std_logic := '0'; 
signal C_49_S_3_L_3_out : std_logic := '0'; 
signal C_49_S_3_L_4_out : std_logic := '0'; 
signal C_49_S_3_L_5_out : std_logic := '0'; 
signal C_49_S_3_L_6_out : std_logic := '0'; 
signal C_49_S_3_L_7_out : std_logic := '0'; 
signal C_49_S_4_L_0_out : std_logic := '0'; 
signal C_49_S_4_L_1_out : std_logic := '0'; 
signal C_49_S_4_L_2_out : std_logic := '0'; 
signal C_49_S_4_L_3_out : std_logic := '0'; 
signal C_49_S_4_L_4_out : std_logic := '0'; 
signal C_49_S_4_L_5_out : std_logic := '0'; 
signal C_49_S_4_L_6_out : std_logic := '0'; 
signal C_49_S_4_L_7_out : std_logic := '0'; 
signal C_50_S_0_L_0_out : std_logic := '0'; 
signal C_50_S_0_L_1_out : std_logic := '0'; 
signal C_50_S_0_L_2_out : std_logic := '0'; 
signal C_50_S_0_L_3_out : std_logic := '0'; 
signal C_50_S_0_L_4_out : std_logic := '0'; 
signal C_50_S_0_L_5_out : std_logic := '0'; 
signal C_50_S_0_L_6_out : std_logic := '0'; 
signal C_50_S_0_L_7_out : std_logic := '0'; 
signal C_50_S_1_L_0_out : std_logic := '0'; 
signal C_50_S_1_L_1_out : std_logic := '0'; 
signal C_50_S_1_L_2_out : std_logic := '0'; 
signal C_50_S_1_L_3_out : std_logic := '0'; 
signal C_50_S_1_L_4_out : std_logic := '0'; 
signal C_50_S_1_L_5_out : std_logic := '0'; 
signal C_50_S_1_L_6_out : std_logic := '0'; 
signal C_50_S_1_L_7_out : std_logic := '0'; 
signal C_50_S_2_L_0_out : std_logic := '0'; 
signal C_50_S_2_L_1_out : std_logic := '0'; 
signal C_50_S_2_L_2_out : std_logic := '0'; 
signal C_50_S_2_L_3_out : std_logic := '0'; 
signal C_50_S_2_L_4_out : std_logic := '0'; 
signal C_50_S_2_L_5_out : std_logic := '0'; 
signal C_50_S_2_L_6_out : std_logic := '0'; 
signal C_50_S_2_L_7_out : std_logic := '0'; 
signal C_50_S_3_L_0_out : std_logic := '0'; 
signal C_50_S_3_L_1_out : std_logic := '0'; 
signal C_50_S_3_L_2_out : std_logic := '0'; 
signal C_50_S_3_L_3_out : std_logic := '0'; 
signal C_50_S_3_L_4_out : std_logic := '0'; 
signal C_50_S_3_L_5_out : std_logic := '0'; 
signal C_50_S_3_L_6_out : std_logic := '0'; 
signal C_50_S_3_L_7_out : std_logic := '0'; 
signal C_50_S_4_L_0_out : std_logic := '0'; 
signal C_50_S_4_L_1_out : std_logic := '0'; 
signal C_50_S_4_L_2_out : std_logic := '0'; 
signal C_50_S_4_L_3_out : std_logic := '0'; 
signal C_50_S_4_L_4_out : std_logic := '0'; 
signal C_50_S_4_L_5_out : std_logic := '0'; 
signal C_50_S_4_L_6_out : std_logic := '0'; 
signal C_50_S_4_L_7_out : std_logic := '0'; 
signal C_51_S_0_L_0_out : std_logic := '0'; 
signal C_51_S_0_L_1_out : std_logic := '0'; 
signal C_51_S_0_L_2_out : std_logic := '0'; 
signal C_51_S_0_L_3_out : std_logic := '0'; 
signal C_51_S_0_L_4_out : std_logic := '0'; 
signal C_51_S_0_L_5_out : std_logic := '0'; 
signal C_51_S_0_L_6_out : std_logic := '0'; 
signal C_51_S_0_L_7_out : std_logic := '0'; 
signal C_51_S_1_L_0_out : std_logic := '0'; 
signal C_51_S_1_L_1_out : std_logic := '0'; 
signal C_51_S_1_L_2_out : std_logic := '0'; 
signal C_51_S_1_L_3_out : std_logic := '0'; 
signal C_51_S_1_L_4_out : std_logic := '0'; 
signal C_51_S_1_L_5_out : std_logic := '0'; 
signal C_51_S_1_L_6_out : std_logic := '0'; 
signal C_51_S_1_L_7_out : std_logic := '0'; 
signal C_51_S_2_L_0_out : std_logic := '0'; 
signal C_51_S_2_L_1_out : std_logic := '0'; 
signal C_51_S_2_L_2_out : std_logic := '0'; 
signal C_51_S_2_L_3_out : std_logic := '0'; 
signal C_51_S_2_L_4_out : std_logic := '0'; 
signal C_51_S_2_L_5_out : std_logic := '0'; 
signal C_51_S_2_L_6_out : std_logic := '0'; 
signal C_51_S_2_L_7_out : std_logic := '0'; 
signal C_51_S_3_L_0_out : std_logic := '0'; 
signal C_51_S_3_L_1_out : std_logic := '0'; 
signal C_51_S_3_L_2_out : std_logic := '0'; 
signal C_51_S_3_L_3_out : std_logic := '0'; 
signal C_51_S_3_L_4_out : std_logic := '0'; 
signal C_51_S_3_L_5_out : std_logic := '0'; 
signal C_51_S_3_L_6_out : std_logic := '0'; 
signal C_51_S_3_L_7_out : std_logic := '0'; 
signal C_51_S_4_L_0_out : std_logic := '0'; 
signal C_51_S_4_L_1_out : std_logic := '0'; 
signal C_51_S_4_L_2_out : std_logic := '0'; 
signal C_51_S_4_L_3_out : std_logic := '0'; 
signal C_51_S_4_L_4_out : std_logic := '0'; 
signal C_51_S_4_L_5_out : std_logic := '0'; 
signal C_51_S_4_L_6_out : std_logic := '0'; 
signal C_51_S_4_L_7_out : std_logic := '0'; 
signal C_52_S_0_L_0_out : std_logic := '0'; 
signal C_52_S_0_L_1_out : std_logic := '0'; 
signal C_52_S_0_L_2_out : std_logic := '0'; 
signal C_52_S_0_L_3_out : std_logic := '0'; 
signal C_52_S_0_L_4_out : std_logic := '0'; 
signal C_52_S_0_L_5_out : std_logic := '0'; 
signal C_52_S_0_L_6_out : std_logic := '0'; 
signal C_52_S_0_L_7_out : std_logic := '0'; 
signal C_52_S_1_L_0_out : std_logic := '0'; 
signal C_52_S_1_L_1_out : std_logic := '0'; 
signal C_52_S_1_L_2_out : std_logic := '0'; 
signal C_52_S_1_L_3_out : std_logic := '0'; 
signal C_52_S_1_L_4_out : std_logic := '0'; 
signal C_52_S_1_L_5_out : std_logic := '0'; 
signal C_52_S_1_L_6_out : std_logic := '0'; 
signal C_52_S_1_L_7_out : std_logic := '0'; 
signal C_52_S_2_L_0_out : std_logic := '0'; 
signal C_52_S_2_L_1_out : std_logic := '0'; 
signal C_52_S_2_L_2_out : std_logic := '0'; 
signal C_52_S_2_L_3_out : std_logic := '0'; 
signal C_52_S_2_L_4_out : std_logic := '0'; 
signal C_52_S_2_L_5_out : std_logic := '0'; 
signal C_52_S_2_L_6_out : std_logic := '0'; 
signal C_52_S_2_L_7_out : std_logic := '0'; 
signal C_52_S_3_L_0_out : std_logic := '0'; 
signal C_52_S_3_L_1_out : std_logic := '0'; 
signal C_52_S_3_L_2_out : std_logic := '0'; 
signal C_52_S_3_L_3_out : std_logic := '0'; 
signal C_52_S_3_L_4_out : std_logic := '0'; 
signal C_52_S_3_L_5_out : std_logic := '0'; 
signal C_52_S_3_L_6_out : std_logic := '0'; 
signal C_52_S_3_L_7_out : std_logic := '0'; 
signal C_52_S_4_L_0_out : std_logic := '0'; 
signal C_52_S_4_L_1_out : std_logic := '0'; 
signal C_52_S_4_L_2_out : std_logic := '0'; 
signal C_52_S_4_L_3_out : std_logic := '0'; 
signal C_52_S_4_L_4_out : std_logic := '0'; 
signal C_52_S_4_L_5_out : std_logic := '0'; 
signal C_52_S_4_L_6_out : std_logic := '0'; 
signal C_52_S_4_L_7_out : std_logic := '0'; 
signal C_53_S_0_L_0_out : std_logic := '0'; 
signal C_53_S_0_L_1_out : std_logic := '0'; 
signal C_53_S_0_L_2_out : std_logic := '0'; 
signal C_53_S_0_L_3_out : std_logic := '0'; 
signal C_53_S_0_L_4_out : std_logic := '0'; 
signal C_53_S_0_L_5_out : std_logic := '0'; 
signal C_53_S_0_L_6_out : std_logic := '0'; 
signal C_53_S_0_L_7_out : std_logic := '0'; 
signal C_53_S_1_L_0_out : std_logic := '0'; 
signal C_53_S_1_L_1_out : std_logic := '0'; 
signal C_53_S_1_L_2_out : std_logic := '0'; 
signal C_53_S_1_L_3_out : std_logic := '0'; 
signal C_53_S_1_L_4_out : std_logic := '0'; 
signal C_53_S_1_L_5_out : std_logic := '0'; 
signal C_53_S_1_L_6_out : std_logic := '0'; 
signal C_53_S_1_L_7_out : std_logic := '0'; 
signal C_53_S_2_L_0_out : std_logic := '0'; 
signal C_53_S_2_L_1_out : std_logic := '0'; 
signal C_53_S_2_L_2_out : std_logic := '0'; 
signal C_53_S_2_L_3_out : std_logic := '0'; 
signal C_53_S_2_L_4_out : std_logic := '0'; 
signal C_53_S_2_L_5_out : std_logic := '0'; 
signal C_53_S_2_L_6_out : std_logic := '0'; 
signal C_53_S_2_L_7_out : std_logic := '0'; 
signal C_53_S_3_L_0_out : std_logic := '0'; 
signal C_53_S_3_L_1_out : std_logic := '0'; 
signal C_53_S_3_L_2_out : std_logic := '0'; 
signal C_53_S_3_L_3_out : std_logic := '0'; 
signal C_53_S_3_L_4_out : std_logic := '0'; 
signal C_53_S_3_L_5_out : std_logic := '0'; 
signal C_53_S_3_L_6_out : std_logic := '0'; 
signal C_53_S_3_L_7_out : std_logic := '0'; 
signal C_53_S_4_L_0_out : std_logic := '0'; 
signal C_53_S_4_L_1_out : std_logic := '0'; 
signal C_53_S_4_L_2_out : std_logic := '0'; 
signal C_53_S_4_L_3_out : std_logic := '0'; 
signal C_53_S_4_L_4_out : std_logic := '0'; 
signal C_53_S_4_L_5_out : std_logic := '0'; 
signal C_53_S_4_L_6_out : std_logic := '0'; 
signal C_53_S_4_L_7_out : std_logic := '0'; 
signal C_54_S_0_L_0_out : std_logic := '0'; 
signal C_54_S_0_L_1_out : std_logic := '0'; 
signal C_54_S_0_L_2_out : std_logic := '0'; 
signal C_54_S_0_L_3_out : std_logic := '0'; 
signal C_54_S_0_L_4_out : std_logic := '0'; 
signal C_54_S_0_L_5_out : std_logic := '0'; 
signal C_54_S_0_L_6_out : std_logic := '0'; 
signal C_54_S_0_L_7_out : std_logic := '0'; 
signal C_54_S_1_L_0_out : std_logic := '0'; 
signal C_54_S_1_L_1_out : std_logic := '0'; 
signal C_54_S_1_L_2_out : std_logic := '0'; 
signal C_54_S_1_L_3_out : std_logic := '0'; 
signal C_54_S_1_L_4_out : std_logic := '0'; 
signal C_54_S_1_L_5_out : std_logic := '0'; 
signal C_54_S_1_L_6_out : std_logic := '0'; 
signal C_54_S_1_L_7_out : std_logic := '0'; 
signal C_54_S_2_L_0_out : std_logic := '0'; 
signal C_54_S_2_L_1_out : std_logic := '0'; 
signal C_54_S_2_L_2_out : std_logic := '0'; 
signal C_54_S_2_L_3_out : std_logic := '0'; 
signal C_54_S_2_L_4_out : std_logic := '0'; 
signal C_54_S_2_L_5_out : std_logic := '0'; 
signal C_54_S_2_L_6_out : std_logic := '0'; 
signal C_54_S_2_L_7_out : std_logic := '0'; 
signal C_54_S_3_L_0_out : std_logic := '0'; 
signal C_54_S_3_L_1_out : std_logic := '0'; 
signal C_54_S_3_L_2_out : std_logic := '0'; 
signal C_54_S_3_L_3_out : std_logic := '0'; 
signal C_54_S_3_L_4_out : std_logic := '0'; 
signal C_54_S_3_L_5_out : std_logic := '0'; 
signal C_54_S_3_L_6_out : std_logic := '0'; 
signal C_54_S_3_L_7_out : std_logic := '0'; 
signal C_54_S_4_L_0_out : std_logic := '0'; 
signal C_54_S_4_L_1_out : std_logic := '0'; 
signal C_54_S_4_L_2_out : std_logic := '0'; 
signal C_54_S_4_L_3_out : std_logic := '0'; 
signal C_54_S_4_L_4_out : std_logic := '0'; 
signal C_54_S_4_L_5_out : std_logic := '0'; 
signal C_54_S_4_L_6_out : std_logic := '0'; 
signal C_54_S_4_L_7_out : std_logic := '0'; 
signal C_55_S_0_L_0_out : std_logic := '0'; 
signal C_55_S_0_L_1_out : std_logic := '0'; 
signal C_55_S_0_L_2_out : std_logic := '0'; 
signal C_55_S_0_L_3_out : std_logic := '0'; 
signal C_55_S_0_L_4_out : std_logic := '0'; 
signal C_55_S_0_L_5_out : std_logic := '0'; 
signal C_55_S_0_L_6_out : std_logic := '0'; 
signal C_55_S_0_L_7_out : std_logic := '0'; 
signal C_55_S_1_L_0_out : std_logic := '0'; 
signal C_55_S_1_L_1_out : std_logic := '0'; 
signal C_55_S_1_L_2_out : std_logic := '0'; 
signal C_55_S_1_L_3_out : std_logic := '0'; 
signal C_55_S_1_L_4_out : std_logic := '0'; 
signal C_55_S_1_L_5_out : std_logic := '0'; 
signal C_55_S_1_L_6_out : std_logic := '0'; 
signal C_55_S_1_L_7_out : std_logic := '0'; 
signal C_55_S_2_L_0_out : std_logic := '0'; 
signal C_55_S_2_L_1_out : std_logic := '0'; 
signal C_55_S_2_L_2_out : std_logic := '0'; 
signal C_55_S_2_L_3_out : std_logic := '0'; 
signal C_55_S_2_L_4_out : std_logic := '0'; 
signal C_55_S_2_L_5_out : std_logic := '0'; 
signal C_55_S_2_L_6_out : std_logic := '0'; 
signal C_55_S_2_L_7_out : std_logic := '0'; 
signal C_55_S_3_L_0_out : std_logic := '0'; 
signal C_55_S_3_L_1_out : std_logic := '0'; 
signal C_55_S_3_L_2_out : std_logic := '0'; 
signal C_55_S_3_L_3_out : std_logic := '0'; 
signal C_55_S_3_L_4_out : std_logic := '0'; 
signal C_55_S_3_L_5_out : std_logic := '0'; 
signal C_55_S_3_L_6_out : std_logic := '0'; 
signal C_55_S_3_L_7_out : std_logic := '0'; 
signal C_55_S_4_L_0_out : std_logic := '0'; 
signal C_55_S_4_L_1_out : std_logic := '0'; 
signal C_55_S_4_L_2_out : std_logic := '0'; 
signal C_55_S_4_L_3_out : std_logic := '0'; 
signal C_55_S_4_L_4_out : std_logic := '0'; 
signal C_55_S_4_L_5_out : std_logic := '0'; 
signal C_55_S_4_L_6_out : std_logic := '0'; 
signal C_55_S_4_L_7_out : std_logic := '0'; 
signal C_56_S_0_L_0_out : std_logic := '0'; 
signal C_56_S_0_L_1_out : std_logic := '0'; 
signal C_56_S_0_L_2_out : std_logic := '0'; 
signal C_56_S_0_L_3_out : std_logic := '0'; 
signal C_56_S_0_L_4_out : std_logic := '0'; 
signal C_56_S_0_L_5_out : std_logic := '0'; 
signal C_56_S_0_L_6_out : std_logic := '0'; 
signal C_56_S_0_L_7_out : std_logic := '0'; 
signal C_56_S_1_L_0_out : std_logic := '0'; 
signal C_56_S_1_L_1_out : std_logic := '0'; 
signal C_56_S_1_L_2_out : std_logic := '0'; 
signal C_56_S_1_L_3_out : std_logic := '0'; 
signal C_56_S_1_L_4_out : std_logic := '0'; 
signal C_56_S_1_L_5_out : std_logic := '0'; 
signal C_56_S_1_L_6_out : std_logic := '0'; 
signal C_56_S_1_L_7_out : std_logic := '0'; 
signal C_56_S_2_L_0_out : std_logic := '0'; 
signal C_56_S_2_L_1_out : std_logic := '0'; 
signal C_56_S_2_L_2_out : std_logic := '0'; 
signal C_56_S_2_L_3_out : std_logic := '0'; 
signal C_56_S_2_L_4_out : std_logic := '0'; 
signal C_56_S_2_L_5_out : std_logic := '0'; 
signal C_56_S_2_L_6_out : std_logic := '0'; 
signal C_56_S_2_L_7_out : std_logic := '0'; 
signal C_56_S_3_L_0_out : std_logic := '0'; 
signal C_56_S_3_L_1_out : std_logic := '0'; 
signal C_56_S_3_L_2_out : std_logic := '0'; 
signal C_56_S_3_L_3_out : std_logic := '0'; 
signal C_56_S_3_L_4_out : std_logic := '0'; 
signal C_56_S_3_L_5_out : std_logic := '0'; 
signal C_56_S_3_L_6_out : std_logic := '0'; 
signal C_56_S_3_L_7_out : std_logic := '0'; 
signal C_56_S_4_L_0_out : std_logic := '0'; 
signal C_56_S_4_L_1_out : std_logic := '0'; 
signal C_56_S_4_L_2_out : std_logic := '0'; 
signal C_56_S_4_L_3_out : std_logic := '0'; 
signal C_56_S_4_L_4_out : std_logic := '0'; 
signal C_56_S_4_L_5_out : std_logic := '0'; 
signal C_56_S_4_L_6_out : std_logic := '0'; 
signal C_56_S_4_L_7_out : std_logic := '0'; 
signal C_57_S_0_L_0_out : std_logic := '0'; 
signal C_57_S_0_L_1_out : std_logic := '0'; 
signal C_57_S_0_L_2_out : std_logic := '0'; 
signal C_57_S_0_L_3_out : std_logic := '0'; 
signal C_57_S_0_L_4_out : std_logic := '0'; 
signal C_57_S_0_L_5_out : std_logic := '0'; 
signal C_57_S_0_L_6_out : std_logic := '0'; 
signal C_57_S_0_L_7_out : std_logic := '0'; 
signal C_57_S_1_L_0_out : std_logic := '0'; 
signal C_57_S_1_L_1_out : std_logic := '0'; 
signal C_57_S_1_L_2_out : std_logic := '0'; 
signal C_57_S_1_L_3_out : std_logic := '0'; 
signal C_57_S_1_L_4_out : std_logic := '0'; 
signal C_57_S_1_L_5_out : std_logic := '0'; 
signal C_57_S_1_L_6_out : std_logic := '0'; 
signal C_57_S_1_L_7_out : std_logic := '0'; 
signal C_57_S_2_L_0_out : std_logic := '0'; 
signal C_57_S_2_L_1_out : std_logic := '0'; 
signal C_57_S_2_L_2_out : std_logic := '0'; 
signal C_57_S_2_L_3_out : std_logic := '0'; 
signal C_57_S_2_L_4_out : std_logic := '0'; 
signal C_57_S_2_L_5_out : std_logic := '0'; 
signal C_57_S_2_L_6_out : std_logic := '0'; 
signal C_57_S_2_L_7_out : std_logic := '0'; 
signal C_57_S_3_L_0_out : std_logic := '0'; 
signal C_57_S_3_L_1_out : std_logic := '0'; 
signal C_57_S_3_L_2_out : std_logic := '0'; 
signal C_57_S_3_L_3_out : std_logic := '0'; 
signal C_57_S_3_L_4_out : std_logic := '0'; 
signal C_57_S_3_L_5_out : std_logic := '0'; 
signal C_57_S_3_L_6_out : std_logic := '0'; 
signal C_57_S_3_L_7_out : std_logic := '0'; 
signal C_57_S_4_L_0_out : std_logic := '0'; 
signal C_57_S_4_L_1_out : std_logic := '0'; 
signal C_57_S_4_L_2_out : std_logic := '0'; 
signal C_57_S_4_L_3_out : std_logic := '0'; 
signal C_57_S_4_L_4_out : std_logic := '0'; 
signal C_57_S_4_L_5_out : std_logic := '0'; 
signal C_57_S_4_L_6_out : std_logic := '0'; 
signal C_57_S_4_L_7_out : std_logic := '0'; 
signal C_58_S_0_L_0_out : std_logic := '0'; 
signal C_58_S_0_L_1_out : std_logic := '0'; 
signal C_58_S_0_L_2_out : std_logic := '0'; 
signal C_58_S_0_L_3_out : std_logic := '0'; 
signal C_58_S_0_L_4_out : std_logic := '0'; 
signal C_58_S_0_L_5_out : std_logic := '0'; 
signal C_58_S_0_L_6_out : std_logic := '0'; 
signal C_58_S_0_L_7_out : std_logic := '0'; 
signal C_58_S_1_L_0_out : std_logic := '0'; 
signal C_58_S_1_L_1_out : std_logic := '0'; 
signal C_58_S_1_L_2_out : std_logic := '0'; 
signal C_58_S_1_L_3_out : std_logic := '0'; 
signal C_58_S_1_L_4_out : std_logic := '0'; 
signal C_58_S_1_L_5_out : std_logic := '0'; 
signal C_58_S_1_L_6_out : std_logic := '0'; 
signal C_58_S_1_L_7_out : std_logic := '0'; 
signal C_58_S_2_L_0_out : std_logic := '0'; 
signal C_58_S_2_L_1_out : std_logic := '0'; 
signal C_58_S_2_L_2_out : std_logic := '0'; 
signal C_58_S_2_L_3_out : std_logic := '0'; 
signal C_58_S_2_L_4_out : std_logic := '0'; 
signal C_58_S_2_L_5_out : std_logic := '0'; 
signal C_58_S_2_L_6_out : std_logic := '0'; 
signal C_58_S_2_L_7_out : std_logic := '0'; 
signal C_58_S_3_L_0_out : std_logic := '0'; 
signal C_58_S_3_L_1_out : std_logic := '0'; 
signal C_58_S_3_L_2_out : std_logic := '0'; 
signal C_58_S_3_L_3_out : std_logic := '0'; 
signal C_58_S_3_L_4_out : std_logic := '0'; 
signal C_58_S_3_L_5_out : std_logic := '0'; 
signal C_58_S_3_L_6_out : std_logic := '0'; 
signal C_58_S_3_L_7_out : std_logic := '0'; 
signal C_58_S_4_L_0_out : std_logic := '0'; 
signal C_58_S_4_L_1_out : std_logic := '0'; 
signal C_58_S_4_L_2_out : std_logic := '0'; 
signal C_58_S_4_L_3_out : std_logic := '0'; 
signal C_58_S_4_L_4_out : std_logic := '0'; 
signal C_58_S_4_L_5_out : std_logic := '0'; 
signal C_58_S_4_L_6_out : std_logic := '0'; 
signal C_58_S_4_L_7_out : std_logic := '0'; 
signal C_59_S_0_L_0_out : std_logic := '0'; 
signal C_59_S_0_L_1_out : std_logic := '0'; 
signal C_59_S_0_L_2_out : std_logic := '0'; 
signal C_59_S_0_L_3_out : std_logic := '0'; 
signal C_59_S_0_L_4_out : std_logic := '0'; 
signal C_59_S_0_L_5_out : std_logic := '0'; 
signal C_59_S_0_L_6_out : std_logic := '0'; 
signal C_59_S_0_L_7_out : std_logic := '0'; 
signal C_59_S_1_L_0_out : std_logic := '0'; 
signal C_59_S_1_L_1_out : std_logic := '0'; 
signal C_59_S_1_L_2_out : std_logic := '0'; 
signal C_59_S_1_L_3_out : std_logic := '0'; 
signal C_59_S_1_L_4_out : std_logic := '0'; 
signal C_59_S_1_L_5_out : std_logic := '0'; 
signal C_59_S_1_L_6_out : std_logic := '0'; 
signal C_59_S_1_L_7_out : std_logic := '0'; 
signal C_59_S_2_L_0_out : std_logic := '0'; 
signal C_59_S_2_L_1_out : std_logic := '0'; 
signal C_59_S_2_L_2_out : std_logic := '0'; 
signal C_59_S_2_L_3_out : std_logic := '0'; 
signal C_59_S_2_L_4_out : std_logic := '0'; 
signal C_59_S_2_L_5_out : std_logic := '0'; 
signal C_59_S_2_L_6_out : std_logic := '0'; 
signal C_59_S_2_L_7_out : std_logic := '0'; 
signal C_59_S_3_L_0_out : std_logic := '0'; 
signal C_59_S_3_L_1_out : std_logic := '0'; 
signal C_59_S_3_L_2_out : std_logic := '0'; 
signal C_59_S_3_L_3_out : std_logic := '0'; 
signal C_59_S_3_L_4_out : std_logic := '0'; 
signal C_59_S_3_L_5_out : std_logic := '0'; 
signal C_59_S_3_L_6_out : std_logic := '0'; 
signal C_59_S_3_L_7_out : std_logic := '0'; 
signal C_59_S_4_L_0_out : std_logic := '0'; 
signal C_59_S_4_L_1_out : std_logic := '0'; 
signal C_59_S_4_L_2_out : std_logic := '0'; 
signal C_59_S_4_L_3_out : std_logic := '0'; 
signal C_59_S_4_L_4_out : std_logic := '0'; 
signal C_59_S_4_L_5_out : std_logic := '0'; 
signal C_59_S_4_L_6_out : std_logic := '0'; 
signal C_59_S_4_L_7_out : std_logic := '0'; 
signal C_60_S_0_L_0_out : std_logic := '0'; 
signal C_60_S_0_L_1_out : std_logic := '0'; 
signal C_60_S_0_L_2_out : std_logic := '0'; 
signal C_60_S_0_L_3_out : std_logic := '0'; 
signal C_60_S_0_L_4_out : std_logic := '0'; 
signal C_60_S_0_L_5_out : std_logic := '0'; 
signal C_60_S_0_L_6_out : std_logic := '0'; 
signal C_60_S_0_L_7_out : std_logic := '0'; 
signal C_60_S_1_L_0_out : std_logic := '0'; 
signal C_60_S_1_L_1_out : std_logic := '0'; 
signal C_60_S_1_L_2_out : std_logic := '0'; 
signal C_60_S_1_L_3_out : std_logic := '0'; 
signal C_60_S_1_L_4_out : std_logic := '0'; 
signal C_60_S_1_L_5_out : std_logic := '0'; 
signal C_60_S_1_L_6_out : std_logic := '0'; 
signal C_60_S_1_L_7_out : std_logic := '0'; 
signal C_60_S_2_L_0_out : std_logic := '0'; 
signal C_60_S_2_L_1_out : std_logic := '0'; 
signal C_60_S_2_L_2_out : std_logic := '0'; 
signal C_60_S_2_L_3_out : std_logic := '0'; 
signal C_60_S_2_L_4_out : std_logic := '0'; 
signal C_60_S_2_L_5_out : std_logic := '0'; 
signal C_60_S_2_L_6_out : std_logic := '0'; 
signal C_60_S_2_L_7_out : std_logic := '0'; 
signal C_60_S_3_L_0_out : std_logic := '0'; 
signal C_60_S_3_L_1_out : std_logic := '0'; 
signal C_60_S_3_L_2_out : std_logic := '0'; 
signal C_60_S_3_L_3_out : std_logic := '0'; 
signal C_60_S_3_L_4_out : std_logic := '0'; 
signal C_60_S_3_L_5_out : std_logic := '0'; 
signal C_60_S_3_L_6_out : std_logic := '0'; 
signal C_60_S_3_L_7_out : std_logic := '0'; 
signal C_60_S_4_L_0_out : std_logic := '0'; 
signal C_60_S_4_L_1_out : std_logic := '0'; 
signal C_60_S_4_L_2_out : std_logic := '0'; 
signal C_60_S_4_L_3_out : std_logic := '0'; 
signal C_60_S_4_L_4_out : std_logic := '0'; 
signal C_60_S_4_L_5_out : std_logic := '0'; 
signal C_60_S_4_L_6_out : std_logic := '0'; 
signal C_60_S_4_L_7_out : std_logic := '0'; 
signal C_61_S_0_L_0_out : std_logic := '0'; 
signal C_61_S_0_L_1_out : std_logic := '0'; 
signal C_61_S_0_L_2_out : std_logic := '0'; 
signal C_61_S_0_L_3_out : std_logic := '0'; 
signal C_61_S_0_L_4_out : std_logic := '0'; 
signal C_61_S_0_L_5_out : std_logic := '0'; 
signal C_61_S_0_L_6_out : std_logic := '0'; 
signal C_61_S_0_L_7_out : std_logic := '0'; 
signal C_61_S_1_L_0_out : std_logic := '0'; 
signal C_61_S_1_L_1_out : std_logic := '0'; 
signal C_61_S_1_L_2_out : std_logic := '0'; 
signal C_61_S_1_L_3_out : std_logic := '0'; 
signal C_61_S_1_L_4_out : std_logic := '0'; 
signal C_61_S_1_L_5_out : std_logic := '0'; 
signal C_61_S_1_L_6_out : std_logic := '0'; 
signal C_61_S_1_L_7_out : std_logic := '0'; 
signal C_61_S_2_L_0_out : std_logic := '0'; 
signal C_61_S_2_L_1_out : std_logic := '0'; 
signal C_61_S_2_L_2_out : std_logic := '0'; 
signal C_61_S_2_L_3_out : std_logic := '0'; 
signal C_61_S_2_L_4_out : std_logic := '0'; 
signal C_61_S_2_L_5_out : std_logic := '0'; 
signal C_61_S_2_L_6_out : std_logic := '0'; 
signal C_61_S_2_L_7_out : std_logic := '0'; 
signal C_61_S_3_L_0_out : std_logic := '0'; 
signal C_61_S_3_L_1_out : std_logic := '0'; 
signal C_61_S_3_L_2_out : std_logic := '0'; 
signal C_61_S_3_L_3_out : std_logic := '0'; 
signal C_61_S_3_L_4_out : std_logic := '0'; 
signal C_61_S_3_L_5_out : std_logic := '0'; 
signal C_61_S_3_L_6_out : std_logic := '0'; 
signal C_61_S_3_L_7_out : std_logic := '0'; 
signal C_61_S_4_L_0_out : std_logic := '0'; 
signal C_61_S_4_L_1_out : std_logic := '0'; 
signal C_61_S_4_L_2_out : std_logic := '0'; 
signal C_61_S_4_L_3_out : std_logic := '0'; 
signal C_61_S_4_L_4_out : std_logic := '0'; 
signal C_61_S_4_L_5_out : std_logic := '0'; 
signal C_61_S_4_L_6_out : std_logic := '0'; 
signal C_61_S_4_L_7_out : std_logic := '0'; 
signal C_62_S_0_L_0_out : std_logic := '0'; 
signal C_62_S_0_L_1_out : std_logic := '0'; 
signal C_62_S_0_L_2_out : std_logic := '0'; 
signal C_62_S_0_L_3_out : std_logic := '0'; 
signal C_62_S_0_L_4_out : std_logic := '0'; 
signal C_62_S_0_L_5_out : std_logic := '0'; 
signal C_62_S_0_L_6_out : std_logic := '0'; 
signal C_62_S_0_L_7_out : std_logic := '0'; 
signal C_62_S_1_L_0_out : std_logic := '0'; 
signal C_62_S_1_L_1_out : std_logic := '0'; 
signal C_62_S_1_L_2_out : std_logic := '0'; 
signal C_62_S_1_L_3_out : std_logic := '0'; 
signal C_62_S_1_L_4_out : std_logic := '0'; 
signal C_62_S_1_L_5_out : std_logic := '0'; 
signal C_62_S_1_L_6_out : std_logic := '0'; 
signal C_62_S_1_L_7_out : std_logic := '0'; 
signal C_62_S_2_L_0_out : std_logic := '0'; 
signal C_62_S_2_L_1_out : std_logic := '0'; 
signal C_62_S_2_L_2_out : std_logic := '0'; 
signal C_62_S_2_L_3_out : std_logic := '0'; 
signal C_62_S_2_L_4_out : std_logic := '0'; 
signal C_62_S_2_L_5_out : std_logic := '0'; 
signal C_62_S_2_L_6_out : std_logic := '0'; 
signal C_62_S_2_L_7_out : std_logic := '0'; 
signal C_62_S_3_L_0_out : std_logic := '0'; 
signal C_62_S_3_L_1_out : std_logic := '0'; 
signal C_62_S_3_L_2_out : std_logic := '0'; 
signal C_62_S_3_L_3_out : std_logic := '0'; 
signal C_62_S_3_L_4_out : std_logic := '0'; 
signal C_62_S_3_L_5_out : std_logic := '0'; 
signal C_62_S_3_L_6_out : std_logic := '0'; 
signal C_62_S_3_L_7_out : std_logic := '0'; 
signal C_62_S_4_L_0_out : std_logic := '0'; 
signal C_62_S_4_L_1_out : std_logic := '0'; 
signal C_62_S_4_L_2_out : std_logic := '0'; 
signal C_62_S_4_L_3_out : std_logic := '0'; 
signal C_62_S_4_L_4_out : std_logic := '0'; 
signal C_62_S_4_L_5_out : std_logic := '0'; 
signal C_62_S_4_L_6_out : std_logic := '0'; 
signal C_62_S_4_L_7_out : std_logic := '0'; 
signal C_63_S_0_L_0_out : std_logic := '0'; 
signal C_63_S_0_L_1_out : std_logic := '0'; 
signal C_63_S_0_L_2_out : std_logic := '0'; 
signal C_63_S_0_L_3_out : std_logic := '0'; 
signal C_63_S_0_L_4_out : std_logic := '0'; 
signal C_63_S_0_L_5_out : std_logic := '0'; 
signal C_63_S_0_L_6_out : std_logic := '0'; 
signal C_63_S_0_L_7_out : std_logic := '0'; 
signal C_63_S_1_L_0_out : std_logic := '0'; 
signal C_63_S_1_L_1_out : std_logic := '0'; 
signal C_63_S_1_L_2_out : std_logic := '0'; 
signal C_63_S_1_L_3_out : std_logic := '0'; 
signal C_63_S_1_L_4_out : std_logic := '0'; 
signal C_63_S_1_L_5_out : std_logic := '0'; 
signal C_63_S_1_L_6_out : std_logic := '0'; 
signal C_63_S_1_L_7_out : std_logic := '0'; 
signal C_63_S_2_L_0_out : std_logic := '0'; 
signal C_63_S_2_L_1_out : std_logic := '0'; 
signal C_63_S_2_L_2_out : std_logic := '0'; 
signal C_63_S_2_L_3_out : std_logic := '0'; 
signal C_63_S_2_L_4_out : std_logic := '0'; 
signal C_63_S_2_L_5_out : std_logic := '0'; 
signal C_63_S_2_L_6_out : std_logic := '0'; 
signal C_63_S_2_L_7_out : std_logic := '0'; 
signal C_63_S_3_L_0_out : std_logic := '0'; 
signal C_63_S_3_L_1_out : std_logic := '0'; 
signal C_63_S_3_L_2_out : std_logic := '0'; 
signal C_63_S_3_L_3_out : std_logic := '0'; 
signal C_63_S_3_L_4_out : std_logic := '0'; 
signal C_63_S_3_L_5_out : std_logic := '0'; 
signal C_63_S_3_L_6_out : std_logic := '0'; 
signal C_63_S_3_L_7_out : std_logic := '0'; 
signal C_63_S_4_L_0_out : std_logic := '0'; 
signal C_63_S_4_L_1_out : std_logic := '0'; 
signal C_63_S_4_L_2_out : std_logic := '0'; 
signal C_63_S_4_L_3_out : std_logic := '0'; 
signal C_63_S_4_L_4_out : std_logic := '0'; 
signal C_63_S_4_L_5_out : std_logic := '0'; 
signal C_63_S_4_L_6_out : std_logic := '0'; 
signal C_63_S_4_L_7_out : std_logic := '0'; 
signal C_64_S_0_L_0_out : std_logic := '0'; 
signal C_64_S_0_L_1_out : std_logic := '0'; 
signal C_64_S_0_L_2_out : std_logic := '0'; 
signal C_64_S_0_L_3_out : std_logic := '0'; 
signal C_64_S_0_L_4_out : std_logic := '0'; 
signal C_64_S_0_L_5_out : std_logic := '0'; 
signal C_64_S_0_L_6_out : std_logic := '0'; 
signal C_64_S_0_L_7_out : std_logic := '0'; 
signal C_64_S_1_L_0_out : std_logic := '0'; 
signal C_64_S_1_L_1_out : std_logic := '0'; 
signal C_64_S_1_L_2_out : std_logic := '0'; 
signal C_64_S_1_L_3_out : std_logic := '0'; 
signal C_64_S_1_L_4_out : std_logic := '0'; 
signal C_64_S_1_L_5_out : std_logic := '0'; 
signal C_64_S_1_L_6_out : std_logic := '0'; 
signal C_64_S_1_L_7_out : std_logic := '0'; 
signal C_64_S_2_L_0_out : std_logic := '0'; 
signal C_64_S_2_L_1_out : std_logic := '0'; 
signal C_64_S_2_L_2_out : std_logic := '0'; 
signal C_64_S_2_L_3_out : std_logic := '0'; 
signal C_64_S_2_L_4_out : std_logic := '0'; 
signal C_64_S_2_L_5_out : std_logic := '0'; 
signal C_64_S_2_L_6_out : std_logic := '0'; 
signal C_64_S_2_L_7_out : std_logic := '0'; 
signal C_64_S_3_L_0_out : std_logic := '0'; 
signal C_64_S_3_L_1_out : std_logic := '0'; 
signal C_64_S_3_L_2_out : std_logic := '0'; 
signal C_64_S_3_L_3_out : std_logic := '0'; 
signal C_64_S_3_L_4_out : std_logic := '0'; 
signal C_64_S_3_L_5_out : std_logic := '0'; 
signal C_64_S_3_L_6_out : std_logic := '0'; 
signal C_64_S_3_L_7_out : std_logic := '0'; 
signal C_64_S_4_L_0_out : std_logic := '0'; 
signal C_64_S_4_L_1_out : std_logic := '0'; 
signal C_64_S_4_L_2_out : std_logic := '0'; 
signal C_64_S_4_L_3_out : std_logic := '0'; 
signal C_64_S_4_L_4_out : std_logic := '0'; 
signal C_64_S_4_L_5_out : std_logic := '0'; 
signal C_64_S_4_L_6_out : std_logic := '0'; 
signal C_64_S_4_L_7_out : std_logic := '0'; 
signal C_65_S_0_L_0_out : std_logic := '0'; 
signal C_65_S_0_L_1_out : std_logic := '0'; 
signal C_65_S_0_L_2_out : std_logic := '0'; 
signal C_65_S_0_L_3_out : std_logic := '0'; 
signal C_65_S_0_L_4_out : std_logic := '0'; 
signal C_65_S_0_L_5_out : std_logic := '0'; 
signal C_65_S_0_L_6_out : std_logic := '0'; 
signal C_65_S_0_L_7_out : std_logic := '0'; 
signal C_65_S_1_L_0_out : std_logic := '0'; 
signal C_65_S_1_L_1_out : std_logic := '0'; 
signal C_65_S_1_L_2_out : std_logic := '0'; 
signal C_65_S_1_L_3_out : std_logic := '0'; 
signal C_65_S_1_L_4_out : std_logic := '0'; 
signal C_65_S_1_L_5_out : std_logic := '0'; 
signal C_65_S_1_L_6_out : std_logic := '0'; 
signal C_65_S_1_L_7_out : std_logic := '0'; 
signal C_65_S_2_L_0_out : std_logic := '0'; 
signal C_65_S_2_L_1_out : std_logic := '0'; 
signal C_65_S_2_L_2_out : std_logic := '0'; 
signal C_65_S_2_L_3_out : std_logic := '0'; 
signal C_65_S_2_L_4_out : std_logic := '0'; 
signal C_65_S_2_L_5_out : std_logic := '0'; 
signal C_65_S_2_L_6_out : std_logic := '0'; 
signal C_65_S_2_L_7_out : std_logic := '0'; 
signal C_65_S_3_L_0_out : std_logic := '0'; 
signal C_65_S_3_L_1_out : std_logic := '0'; 
signal C_65_S_3_L_2_out : std_logic := '0'; 
signal C_65_S_3_L_3_out : std_logic := '0'; 
signal C_65_S_3_L_4_out : std_logic := '0'; 
signal C_65_S_3_L_5_out : std_logic := '0'; 
signal C_65_S_3_L_6_out : std_logic := '0'; 
signal C_65_S_3_L_7_out : std_logic := '0'; 
signal C_65_S_4_L_0_out : std_logic := '0'; 
signal C_65_S_4_L_1_out : std_logic := '0'; 
signal C_65_S_4_L_2_out : std_logic := '0'; 
signal C_65_S_4_L_3_out : std_logic := '0'; 
signal C_65_S_4_L_4_out : std_logic := '0'; 
signal C_65_S_4_L_5_out : std_logic := '0'; 
signal C_65_S_4_L_6_out : std_logic := '0'; 
signal C_65_S_4_L_7_out : std_logic := '0'; 
signal C_66_S_0_L_0_out : std_logic := '0'; 
signal C_66_S_0_L_1_out : std_logic := '0'; 
signal C_66_S_0_L_2_out : std_logic := '0'; 
signal C_66_S_0_L_3_out : std_logic := '0'; 
signal C_66_S_0_L_4_out : std_logic := '0'; 
signal C_66_S_0_L_5_out : std_logic := '0'; 
signal C_66_S_0_L_6_out : std_logic := '0'; 
signal C_66_S_0_L_7_out : std_logic := '0'; 
signal C_66_S_1_L_0_out : std_logic := '0'; 
signal C_66_S_1_L_1_out : std_logic := '0'; 
signal C_66_S_1_L_2_out : std_logic := '0'; 
signal C_66_S_1_L_3_out : std_logic := '0'; 
signal C_66_S_1_L_4_out : std_logic := '0'; 
signal C_66_S_1_L_5_out : std_logic := '0'; 
signal C_66_S_1_L_6_out : std_logic := '0'; 
signal C_66_S_1_L_7_out : std_logic := '0'; 
signal C_66_S_2_L_0_out : std_logic := '0'; 
signal C_66_S_2_L_1_out : std_logic := '0'; 
signal C_66_S_2_L_2_out : std_logic := '0'; 
signal C_66_S_2_L_3_out : std_logic := '0'; 
signal C_66_S_2_L_4_out : std_logic := '0'; 
signal C_66_S_2_L_5_out : std_logic := '0'; 
signal C_66_S_2_L_6_out : std_logic := '0'; 
signal C_66_S_2_L_7_out : std_logic := '0'; 
signal C_66_S_3_L_0_out : std_logic := '0'; 
signal C_66_S_3_L_1_out : std_logic := '0'; 
signal C_66_S_3_L_2_out : std_logic := '0'; 
signal C_66_S_3_L_3_out : std_logic := '0'; 
signal C_66_S_3_L_4_out : std_logic := '0'; 
signal C_66_S_3_L_5_out : std_logic := '0'; 
signal C_66_S_3_L_6_out : std_logic := '0'; 
signal C_66_S_3_L_7_out : std_logic := '0'; 
signal C_66_S_4_L_0_out : std_logic := '0'; 
signal C_66_S_4_L_1_out : std_logic := '0'; 
signal C_66_S_4_L_2_out : std_logic := '0'; 
signal C_66_S_4_L_3_out : std_logic := '0'; 
signal C_66_S_4_L_4_out : std_logic := '0'; 
signal C_66_S_4_L_5_out : std_logic := '0'; 
signal C_66_S_4_L_6_out : std_logic := '0'; 
signal C_66_S_4_L_7_out : std_logic := '0'; 
signal C_67_S_0_L_0_out : std_logic := '0'; 
signal C_67_S_0_L_1_out : std_logic := '0'; 
signal C_67_S_0_L_2_out : std_logic := '0'; 
signal C_67_S_0_L_3_out : std_logic := '0'; 
signal C_67_S_0_L_4_out : std_logic := '0'; 
signal C_67_S_0_L_5_out : std_logic := '0'; 
signal C_67_S_0_L_6_out : std_logic := '0'; 
signal C_67_S_0_L_7_out : std_logic := '0'; 
signal C_67_S_1_L_0_out : std_logic := '0'; 
signal C_67_S_1_L_1_out : std_logic := '0'; 
signal C_67_S_1_L_2_out : std_logic := '0'; 
signal C_67_S_1_L_3_out : std_logic := '0'; 
signal C_67_S_1_L_4_out : std_logic := '0'; 
signal C_67_S_1_L_5_out : std_logic := '0'; 
signal C_67_S_1_L_6_out : std_logic := '0'; 
signal C_67_S_1_L_7_out : std_logic := '0'; 
signal C_67_S_2_L_0_out : std_logic := '0'; 
signal C_67_S_2_L_1_out : std_logic := '0'; 
signal C_67_S_2_L_2_out : std_logic := '0'; 
signal C_67_S_2_L_3_out : std_logic := '0'; 
signal C_67_S_2_L_4_out : std_logic := '0'; 
signal C_67_S_2_L_5_out : std_logic := '0'; 
signal C_67_S_2_L_6_out : std_logic := '0'; 
signal C_67_S_2_L_7_out : std_logic := '0'; 
signal C_67_S_3_L_0_out : std_logic := '0'; 
signal C_67_S_3_L_1_out : std_logic := '0'; 
signal C_67_S_3_L_2_out : std_logic := '0'; 
signal C_67_S_3_L_3_out : std_logic := '0'; 
signal C_67_S_3_L_4_out : std_logic := '0'; 
signal C_67_S_3_L_5_out : std_logic := '0'; 
signal C_67_S_3_L_6_out : std_logic := '0'; 
signal C_67_S_3_L_7_out : std_logic := '0'; 
signal C_67_S_4_L_0_out : std_logic := '0'; 
signal C_67_S_4_L_1_out : std_logic := '0'; 
signal C_67_S_4_L_2_out : std_logic := '0'; 
signal C_67_S_4_L_3_out : std_logic := '0'; 
signal C_67_S_4_L_4_out : std_logic := '0'; 
signal C_67_S_4_L_5_out : std_logic := '0'; 
signal C_67_S_4_L_6_out : std_logic := '0'; 
signal C_67_S_4_L_7_out : std_logic := '0'; 
signal C_68_S_0_L_0_out : std_logic := '0'; 
signal C_68_S_0_L_1_out : std_logic := '0'; 
signal C_68_S_0_L_2_out : std_logic := '0'; 
signal C_68_S_0_L_3_out : std_logic := '0'; 
signal C_68_S_0_L_4_out : std_logic := '0'; 
signal C_68_S_0_L_5_out : std_logic := '0'; 
signal C_68_S_0_L_6_out : std_logic := '0'; 
signal C_68_S_0_L_7_out : std_logic := '0'; 
signal C_68_S_1_L_0_out : std_logic := '0'; 
signal C_68_S_1_L_1_out : std_logic := '0'; 
signal C_68_S_1_L_2_out : std_logic := '0'; 
signal C_68_S_1_L_3_out : std_logic := '0'; 
signal C_68_S_1_L_4_out : std_logic := '0'; 
signal C_68_S_1_L_5_out : std_logic := '0'; 
signal C_68_S_1_L_6_out : std_logic := '0'; 
signal C_68_S_1_L_7_out : std_logic := '0'; 
signal C_68_S_2_L_0_out : std_logic := '0'; 
signal C_68_S_2_L_1_out : std_logic := '0'; 
signal C_68_S_2_L_2_out : std_logic := '0'; 
signal C_68_S_2_L_3_out : std_logic := '0'; 
signal C_68_S_2_L_4_out : std_logic := '0'; 
signal C_68_S_2_L_5_out : std_logic := '0'; 
signal C_68_S_2_L_6_out : std_logic := '0'; 
signal C_68_S_2_L_7_out : std_logic := '0'; 
signal C_68_S_3_L_0_out : std_logic := '0'; 
signal C_68_S_3_L_1_out : std_logic := '0'; 
signal C_68_S_3_L_2_out : std_logic := '0'; 
signal C_68_S_3_L_3_out : std_logic := '0'; 
signal C_68_S_3_L_4_out : std_logic := '0'; 
signal C_68_S_3_L_5_out : std_logic := '0'; 
signal C_68_S_3_L_6_out : std_logic := '0'; 
signal C_68_S_3_L_7_out : std_logic := '0'; 
signal C_68_S_4_L_0_out : std_logic := '0'; 
signal C_68_S_4_L_1_out : std_logic := '0'; 
signal C_68_S_4_L_2_out : std_logic := '0'; 
signal C_68_S_4_L_3_out : std_logic := '0'; 
signal C_68_S_4_L_4_out : std_logic := '0'; 
signal C_68_S_4_L_5_out : std_logic := '0'; 
signal C_68_S_4_L_6_out : std_logic := '0'; 
signal C_68_S_4_L_7_out : std_logic := '0'; 
signal C_69_S_0_L_0_out : std_logic := '0'; 
signal C_69_S_0_L_1_out : std_logic := '0'; 
signal C_69_S_0_L_2_out : std_logic := '0'; 
signal C_69_S_0_L_3_out : std_logic := '0'; 
signal C_69_S_0_L_4_out : std_logic := '0'; 
signal C_69_S_0_L_5_out : std_logic := '0'; 
signal C_69_S_0_L_6_out : std_logic := '0'; 
signal C_69_S_0_L_7_out : std_logic := '0'; 
signal C_69_S_1_L_0_out : std_logic := '0'; 
signal C_69_S_1_L_1_out : std_logic := '0'; 
signal C_69_S_1_L_2_out : std_logic := '0'; 
signal C_69_S_1_L_3_out : std_logic := '0'; 
signal C_69_S_1_L_4_out : std_logic := '0'; 
signal C_69_S_1_L_5_out : std_logic := '0'; 
signal C_69_S_1_L_6_out : std_logic := '0'; 
signal C_69_S_1_L_7_out : std_logic := '0'; 
signal C_69_S_2_L_0_out : std_logic := '0'; 
signal C_69_S_2_L_1_out : std_logic := '0'; 
signal C_69_S_2_L_2_out : std_logic := '0'; 
signal C_69_S_2_L_3_out : std_logic := '0'; 
signal C_69_S_2_L_4_out : std_logic := '0'; 
signal C_69_S_2_L_5_out : std_logic := '0'; 
signal C_69_S_2_L_6_out : std_logic := '0'; 
signal C_69_S_2_L_7_out : std_logic := '0'; 
signal C_69_S_3_L_0_out : std_logic := '0'; 
signal C_69_S_3_L_1_out : std_logic := '0'; 
signal C_69_S_3_L_2_out : std_logic := '0'; 
signal C_69_S_3_L_3_out : std_logic := '0'; 
signal C_69_S_3_L_4_out : std_logic := '0'; 
signal C_69_S_3_L_5_out : std_logic := '0'; 
signal C_69_S_3_L_6_out : std_logic := '0'; 
signal C_69_S_3_L_7_out : std_logic := '0'; 
signal C_69_S_4_L_0_out : std_logic := '0'; 
signal C_69_S_4_L_1_out : std_logic := '0'; 
signal C_69_S_4_L_2_out : std_logic := '0'; 
signal C_69_S_4_L_3_out : std_logic := '0'; 
signal C_69_S_4_L_4_out : std_logic := '0'; 
signal C_69_S_4_L_5_out : std_logic := '0'; 
signal C_69_S_4_L_6_out : std_logic := '0'; 
signal C_69_S_4_L_7_out : std_logic := '0'; 
signal C_70_S_0_L_0_out : std_logic := '0'; 
signal C_70_S_0_L_1_out : std_logic := '0'; 
signal C_70_S_0_L_2_out : std_logic := '0'; 
signal C_70_S_0_L_3_out : std_logic := '0'; 
signal C_70_S_0_L_4_out : std_logic := '0'; 
signal C_70_S_0_L_5_out : std_logic := '0'; 
signal C_70_S_0_L_6_out : std_logic := '0'; 
signal C_70_S_0_L_7_out : std_logic := '0'; 
signal C_70_S_1_L_0_out : std_logic := '0'; 
signal C_70_S_1_L_1_out : std_logic := '0'; 
signal C_70_S_1_L_2_out : std_logic := '0'; 
signal C_70_S_1_L_3_out : std_logic := '0'; 
signal C_70_S_1_L_4_out : std_logic := '0'; 
signal C_70_S_1_L_5_out : std_logic := '0'; 
signal C_70_S_1_L_6_out : std_logic := '0'; 
signal C_70_S_1_L_7_out : std_logic := '0'; 
signal C_70_S_2_L_0_out : std_logic := '0'; 
signal C_70_S_2_L_1_out : std_logic := '0'; 
signal C_70_S_2_L_2_out : std_logic := '0'; 
signal C_70_S_2_L_3_out : std_logic := '0'; 
signal C_70_S_2_L_4_out : std_logic := '0'; 
signal C_70_S_2_L_5_out : std_logic := '0'; 
signal C_70_S_2_L_6_out : std_logic := '0'; 
signal C_70_S_2_L_7_out : std_logic := '0'; 
signal C_70_S_3_L_0_out : std_logic := '0'; 
signal C_70_S_3_L_1_out : std_logic := '0'; 
signal C_70_S_3_L_2_out : std_logic := '0'; 
signal C_70_S_3_L_3_out : std_logic := '0'; 
signal C_70_S_3_L_4_out : std_logic := '0'; 
signal C_70_S_3_L_5_out : std_logic := '0'; 
signal C_70_S_3_L_6_out : std_logic := '0'; 
signal C_70_S_3_L_7_out : std_logic := '0'; 
signal C_70_S_4_L_0_out : std_logic := '0'; 
signal C_70_S_4_L_1_out : std_logic := '0'; 
signal C_70_S_4_L_2_out : std_logic := '0'; 
signal C_70_S_4_L_3_out : std_logic := '0'; 
signal C_70_S_4_L_4_out : std_logic := '0'; 
signal C_70_S_4_L_5_out : std_logic := '0'; 
signal C_70_S_4_L_6_out : std_logic := '0'; 
signal C_70_S_4_L_7_out : std_logic := '0'; 
signal C_71_S_0_L_0_out : std_logic := '0'; 
signal C_71_S_0_L_1_out : std_logic := '0'; 
signal C_71_S_0_L_2_out : std_logic := '0'; 
signal C_71_S_0_L_3_out : std_logic := '0'; 
signal C_71_S_0_L_4_out : std_logic := '0'; 
signal C_71_S_0_L_5_out : std_logic := '0'; 
signal C_71_S_0_L_6_out : std_logic := '0'; 
signal C_71_S_0_L_7_out : std_logic := '0'; 
signal C_71_S_1_L_0_out : std_logic := '0'; 
signal C_71_S_1_L_1_out : std_logic := '0'; 
signal C_71_S_1_L_2_out : std_logic := '0'; 
signal C_71_S_1_L_3_out : std_logic := '0'; 
signal C_71_S_1_L_4_out : std_logic := '0'; 
signal C_71_S_1_L_5_out : std_logic := '0'; 
signal C_71_S_1_L_6_out : std_logic := '0'; 
signal C_71_S_1_L_7_out : std_logic := '0'; 
signal C_71_S_2_L_0_out : std_logic := '0'; 
signal C_71_S_2_L_1_out : std_logic := '0'; 
signal C_71_S_2_L_2_out : std_logic := '0'; 
signal C_71_S_2_L_3_out : std_logic := '0'; 
signal C_71_S_2_L_4_out : std_logic := '0'; 
signal C_71_S_2_L_5_out : std_logic := '0'; 
signal C_71_S_2_L_6_out : std_logic := '0'; 
signal C_71_S_2_L_7_out : std_logic := '0'; 
signal C_71_S_3_L_0_out : std_logic := '0'; 
signal C_71_S_3_L_1_out : std_logic := '0'; 
signal C_71_S_3_L_2_out : std_logic := '0'; 
signal C_71_S_3_L_3_out : std_logic := '0'; 
signal C_71_S_3_L_4_out : std_logic := '0'; 
signal C_71_S_3_L_5_out : std_logic := '0'; 
signal C_71_S_3_L_6_out : std_logic := '0'; 
signal C_71_S_3_L_7_out : std_logic := '0'; 
signal C_71_S_4_L_0_out : std_logic := '0'; 
signal C_71_S_4_L_1_out : std_logic := '0'; 
signal C_71_S_4_L_2_out : std_logic := '0'; 
signal C_71_S_4_L_3_out : std_logic := '0'; 
signal C_71_S_4_L_4_out : std_logic := '0'; 
signal C_71_S_4_L_5_out : std_logic := '0'; 
signal C_71_S_4_L_6_out : std_logic := '0'; 
signal C_71_S_4_L_7_out : std_logic := '0'; 
signal C_72_S_0_L_0_out : std_logic := '0'; 
signal C_72_S_0_L_1_out : std_logic := '0'; 
signal C_72_S_0_L_2_out : std_logic := '0'; 
signal C_72_S_0_L_3_out : std_logic := '0'; 
signal C_72_S_0_L_4_out : std_logic := '0'; 
signal C_72_S_0_L_5_out : std_logic := '0'; 
signal C_72_S_0_L_6_out : std_logic := '0'; 
signal C_72_S_0_L_7_out : std_logic := '0'; 
signal C_72_S_1_L_0_out : std_logic := '0'; 
signal C_72_S_1_L_1_out : std_logic := '0'; 
signal C_72_S_1_L_2_out : std_logic := '0'; 
signal C_72_S_1_L_3_out : std_logic := '0'; 
signal C_72_S_1_L_4_out : std_logic := '0'; 
signal C_72_S_1_L_5_out : std_logic := '0'; 
signal C_72_S_1_L_6_out : std_logic := '0'; 
signal C_72_S_1_L_7_out : std_logic := '0'; 
signal C_72_S_2_L_0_out : std_logic := '0'; 
signal C_72_S_2_L_1_out : std_logic := '0'; 
signal C_72_S_2_L_2_out : std_logic := '0'; 
signal C_72_S_2_L_3_out : std_logic := '0'; 
signal C_72_S_2_L_4_out : std_logic := '0'; 
signal C_72_S_2_L_5_out : std_logic := '0'; 
signal C_72_S_2_L_6_out : std_logic := '0'; 
signal C_72_S_2_L_7_out : std_logic := '0'; 
signal C_72_S_3_L_0_out : std_logic := '0'; 
signal C_72_S_3_L_1_out : std_logic := '0'; 
signal C_72_S_3_L_2_out : std_logic := '0'; 
signal C_72_S_3_L_3_out : std_logic := '0'; 
signal C_72_S_3_L_4_out : std_logic := '0'; 
signal C_72_S_3_L_5_out : std_logic := '0'; 
signal C_72_S_3_L_6_out : std_logic := '0'; 
signal C_72_S_3_L_7_out : std_logic := '0'; 
signal C_72_S_4_L_0_out : std_logic := '0'; 
signal C_72_S_4_L_1_out : std_logic := '0'; 
signal C_72_S_4_L_2_out : std_logic := '0'; 
signal C_72_S_4_L_3_out : std_logic := '0'; 
signal C_72_S_4_L_4_out : std_logic := '0'; 
signal C_72_S_4_L_5_out : std_logic := '0'; 
signal C_72_S_4_L_6_out : std_logic := '0'; 
signal C_72_S_4_L_7_out : std_logic := '0'; 
signal C_73_S_0_L_0_out : std_logic := '0'; 
signal C_73_S_0_L_1_out : std_logic := '0'; 
signal C_73_S_0_L_2_out : std_logic := '0'; 
signal C_73_S_0_L_3_out : std_logic := '0'; 
signal C_73_S_0_L_4_out : std_logic := '0'; 
signal C_73_S_0_L_5_out : std_logic := '0'; 
signal C_73_S_0_L_6_out : std_logic := '0'; 
signal C_73_S_0_L_7_out : std_logic := '0'; 
signal C_73_S_1_L_0_out : std_logic := '0'; 
signal C_73_S_1_L_1_out : std_logic := '0'; 
signal C_73_S_1_L_2_out : std_logic := '0'; 
signal C_73_S_1_L_3_out : std_logic := '0'; 
signal C_73_S_1_L_4_out : std_logic := '0'; 
signal C_73_S_1_L_5_out : std_logic := '0'; 
signal C_73_S_1_L_6_out : std_logic := '0'; 
signal C_73_S_1_L_7_out : std_logic := '0'; 
signal C_73_S_2_L_0_out : std_logic := '0'; 
signal C_73_S_2_L_1_out : std_logic := '0'; 
signal C_73_S_2_L_2_out : std_logic := '0'; 
signal C_73_S_2_L_3_out : std_logic := '0'; 
signal C_73_S_2_L_4_out : std_logic := '0'; 
signal C_73_S_2_L_5_out : std_logic := '0'; 
signal C_73_S_2_L_6_out : std_logic := '0'; 
signal C_73_S_2_L_7_out : std_logic := '0'; 
signal C_73_S_3_L_0_out : std_logic := '0'; 
signal C_73_S_3_L_1_out : std_logic := '0'; 
signal C_73_S_3_L_2_out : std_logic := '0'; 
signal C_73_S_3_L_3_out : std_logic := '0'; 
signal C_73_S_3_L_4_out : std_logic := '0'; 
signal C_73_S_3_L_5_out : std_logic := '0'; 
signal C_73_S_3_L_6_out : std_logic := '0'; 
signal C_73_S_3_L_7_out : std_logic := '0'; 
signal C_73_S_4_L_0_out : std_logic := '0'; 
signal C_73_S_4_L_1_out : std_logic := '0'; 
signal C_73_S_4_L_2_out : std_logic := '0'; 
signal C_73_S_4_L_3_out : std_logic := '0'; 
signal C_73_S_4_L_4_out : std_logic := '0'; 
signal C_73_S_4_L_5_out : std_logic := '0'; 
signal C_73_S_4_L_6_out : std_logic := '0'; 
signal C_73_S_4_L_7_out : std_logic := '0'; 
signal C_74_S_0_L_0_out : std_logic := '0'; 
signal C_74_S_0_L_1_out : std_logic := '0'; 
signal C_74_S_0_L_2_out : std_logic := '0'; 
signal C_74_S_0_L_3_out : std_logic := '0'; 
signal C_74_S_0_L_4_out : std_logic := '0'; 
signal C_74_S_0_L_5_out : std_logic := '0'; 
signal C_74_S_0_L_6_out : std_logic := '0'; 
signal C_74_S_0_L_7_out : std_logic := '0'; 
signal C_74_S_1_L_0_out : std_logic := '0'; 
signal C_74_S_1_L_1_out : std_logic := '0'; 
signal C_74_S_1_L_2_out : std_logic := '0'; 
signal C_74_S_1_L_3_out : std_logic := '0'; 
signal C_74_S_1_L_4_out : std_logic := '0'; 
signal C_74_S_1_L_5_out : std_logic := '0'; 
signal C_74_S_1_L_6_out : std_logic := '0'; 
signal C_74_S_1_L_7_out : std_logic := '0'; 
signal C_74_S_2_L_0_out : std_logic := '0'; 
signal C_74_S_2_L_1_out : std_logic := '0'; 
signal C_74_S_2_L_2_out : std_logic := '0'; 
signal C_74_S_2_L_3_out : std_logic := '0'; 
signal C_74_S_2_L_4_out : std_logic := '0'; 
signal C_74_S_2_L_5_out : std_logic := '0'; 
signal C_74_S_2_L_6_out : std_logic := '0'; 
signal C_74_S_2_L_7_out : std_logic := '0'; 
signal C_74_S_3_L_0_out : std_logic := '0'; 
signal C_74_S_3_L_1_out : std_logic := '0'; 
signal C_74_S_3_L_2_out : std_logic := '0'; 
signal C_74_S_3_L_3_out : std_logic := '0'; 
signal C_74_S_3_L_4_out : std_logic := '0'; 
signal C_74_S_3_L_5_out : std_logic := '0'; 
signal C_74_S_3_L_6_out : std_logic := '0'; 
signal C_74_S_3_L_7_out : std_logic := '0'; 
signal C_74_S_4_L_0_out : std_logic := '0'; 
signal C_74_S_4_L_1_out : std_logic := '0'; 
signal C_74_S_4_L_2_out : std_logic := '0'; 
signal C_74_S_4_L_3_out : std_logic := '0'; 
signal C_74_S_4_L_4_out : std_logic := '0'; 
signal C_74_S_4_L_5_out : std_logic := '0'; 
signal C_74_S_4_L_6_out : std_logic := '0'; 
signal C_74_S_4_L_7_out : std_logic := '0'; 
signal C_75_S_0_L_0_out : std_logic := '0'; 
signal C_75_S_0_L_1_out : std_logic := '0'; 
signal C_75_S_0_L_2_out : std_logic := '0'; 
signal C_75_S_0_L_3_out : std_logic := '0'; 
signal C_75_S_0_L_4_out : std_logic := '0'; 
signal C_75_S_0_L_5_out : std_logic := '0'; 
signal C_75_S_0_L_6_out : std_logic := '0'; 
signal C_75_S_0_L_7_out : std_logic := '0'; 
signal C_75_S_1_L_0_out : std_logic := '0'; 
signal C_75_S_1_L_1_out : std_logic := '0'; 
signal C_75_S_1_L_2_out : std_logic := '0'; 
signal C_75_S_1_L_3_out : std_logic := '0'; 
signal C_75_S_1_L_4_out : std_logic := '0'; 
signal C_75_S_1_L_5_out : std_logic := '0'; 
signal C_75_S_1_L_6_out : std_logic := '0'; 
signal C_75_S_1_L_7_out : std_logic := '0'; 
signal C_75_S_2_L_0_out : std_logic := '0'; 
signal C_75_S_2_L_1_out : std_logic := '0'; 
signal C_75_S_2_L_2_out : std_logic := '0'; 
signal C_75_S_2_L_3_out : std_logic := '0'; 
signal C_75_S_2_L_4_out : std_logic := '0'; 
signal C_75_S_2_L_5_out : std_logic := '0'; 
signal C_75_S_2_L_6_out : std_logic := '0'; 
signal C_75_S_2_L_7_out : std_logic := '0'; 
signal C_75_S_3_L_0_out : std_logic := '0'; 
signal C_75_S_3_L_1_out : std_logic := '0'; 
signal C_75_S_3_L_2_out : std_logic := '0'; 
signal C_75_S_3_L_3_out : std_logic := '0'; 
signal C_75_S_3_L_4_out : std_logic := '0'; 
signal C_75_S_3_L_5_out : std_logic := '0'; 
signal C_75_S_3_L_6_out : std_logic := '0'; 
signal C_75_S_3_L_7_out : std_logic := '0'; 
signal C_75_S_4_L_0_out : std_logic := '0'; 
signal C_75_S_4_L_1_out : std_logic := '0'; 
signal C_75_S_4_L_2_out : std_logic := '0'; 
signal C_75_S_4_L_3_out : std_logic := '0'; 
signal C_75_S_4_L_4_out : std_logic := '0'; 
signal C_75_S_4_L_5_out : std_logic := '0'; 
signal C_75_S_4_L_6_out : std_logic := '0'; 
signal C_75_S_4_L_7_out : std_logic := '0'; 
signal C_76_S_0_L_0_out : std_logic := '0'; 
signal C_76_S_0_L_1_out : std_logic := '0'; 
signal C_76_S_0_L_2_out : std_logic := '0'; 
signal C_76_S_0_L_3_out : std_logic := '0'; 
signal C_76_S_0_L_4_out : std_logic := '0'; 
signal C_76_S_0_L_5_out : std_logic := '0'; 
signal C_76_S_0_L_6_out : std_logic := '0'; 
signal C_76_S_0_L_7_out : std_logic := '0'; 
signal C_76_S_1_L_0_out : std_logic := '0'; 
signal C_76_S_1_L_1_out : std_logic := '0'; 
signal C_76_S_1_L_2_out : std_logic := '0'; 
signal C_76_S_1_L_3_out : std_logic := '0'; 
signal C_76_S_1_L_4_out : std_logic := '0'; 
signal C_76_S_1_L_5_out : std_logic := '0'; 
signal C_76_S_1_L_6_out : std_logic := '0'; 
signal C_76_S_1_L_7_out : std_logic := '0'; 
signal C_76_S_2_L_0_out : std_logic := '0'; 
signal C_76_S_2_L_1_out : std_logic := '0'; 
signal C_76_S_2_L_2_out : std_logic := '0'; 
signal C_76_S_2_L_3_out : std_logic := '0'; 
signal C_76_S_2_L_4_out : std_logic := '0'; 
signal C_76_S_2_L_5_out : std_logic := '0'; 
signal C_76_S_2_L_6_out : std_logic := '0'; 
signal C_76_S_2_L_7_out : std_logic := '0'; 
signal C_76_S_3_L_0_out : std_logic := '0'; 
signal C_76_S_3_L_1_out : std_logic := '0'; 
signal C_76_S_3_L_2_out : std_logic := '0'; 
signal C_76_S_3_L_3_out : std_logic := '0'; 
signal C_76_S_3_L_4_out : std_logic := '0'; 
signal C_76_S_3_L_5_out : std_logic := '0'; 
signal C_76_S_3_L_6_out : std_logic := '0'; 
signal C_76_S_3_L_7_out : std_logic := '0'; 
signal C_76_S_4_L_0_out : std_logic := '0'; 
signal C_76_S_4_L_1_out : std_logic := '0'; 
signal C_76_S_4_L_2_out : std_logic := '0'; 
signal C_76_S_4_L_3_out : std_logic := '0'; 
signal C_76_S_4_L_4_out : std_logic := '0'; 
signal C_76_S_4_L_5_out : std_logic := '0'; 
signal C_76_S_4_L_6_out : std_logic := '0'; 
signal C_76_S_4_L_7_out : std_logic := '0'; 
signal C_77_S_0_L_0_out : std_logic := '0'; 
signal C_77_S_0_L_1_out : std_logic := '0'; 
signal C_77_S_0_L_2_out : std_logic := '0'; 
signal C_77_S_0_L_3_out : std_logic := '0'; 
signal C_77_S_0_L_4_out : std_logic := '0'; 
signal C_77_S_0_L_5_out : std_logic := '0'; 
signal C_77_S_0_L_6_out : std_logic := '0'; 
signal C_77_S_0_L_7_out : std_logic := '0'; 
signal C_77_S_1_L_0_out : std_logic := '0'; 
signal C_77_S_1_L_1_out : std_logic := '0'; 
signal C_77_S_1_L_2_out : std_logic := '0'; 
signal C_77_S_1_L_3_out : std_logic := '0'; 
signal C_77_S_1_L_4_out : std_logic := '0'; 
signal C_77_S_1_L_5_out : std_logic := '0'; 
signal C_77_S_1_L_6_out : std_logic := '0'; 
signal C_77_S_1_L_7_out : std_logic := '0'; 
signal C_77_S_2_L_0_out : std_logic := '0'; 
signal C_77_S_2_L_1_out : std_logic := '0'; 
signal C_77_S_2_L_2_out : std_logic := '0'; 
signal C_77_S_2_L_3_out : std_logic := '0'; 
signal C_77_S_2_L_4_out : std_logic := '0'; 
signal C_77_S_2_L_5_out : std_logic := '0'; 
signal C_77_S_2_L_6_out : std_logic := '0'; 
signal C_77_S_2_L_7_out : std_logic := '0'; 
signal C_77_S_3_L_0_out : std_logic := '0'; 
signal C_77_S_3_L_1_out : std_logic := '0'; 
signal C_77_S_3_L_2_out : std_logic := '0'; 
signal C_77_S_3_L_3_out : std_logic := '0'; 
signal C_77_S_3_L_4_out : std_logic := '0'; 
signal C_77_S_3_L_5_out : std_logic := '0'; 
signal C_77_S_3_L_6_out : std_logic := '0'; 
signal C_77_S_3_L_7_out : std_logic := '0'; 
signal C_77_S_4_L_0_out : std_logic := '0'; 
signal C_77_S_4_L_1_out : std_logic := '0'; 
signal C_77_S_4_L_2_out : std_logic := '0'; 
signal C_77_S_4_L_3_out : std_logic := '0'; 
signal C_77_S_4_L_4_out : std_logic := '0'; 
signal C_77_S_4_L_5_out : std_logic := '0'; 
signal C_77_S_4_L_6_out : std_logic := '0'; 
signal C_77_S_4_L_7_out : std_logic := '0'; 
signal C_78_S_0_L_0_out : std_logic := '0'; 
signal C_78_S_0_L_1_out : std_logic := '0'; 
signal C_78_S_0_L_2_out : std_logic := '0'; 
signal C_78_S_0_L_3_out : std_logic := '0'; 
signal C_78_S_0_L_4_out : std_logic := '0'; 
signal C_78_S_0_L_5_out : std_logic := '0'; 
signal C_78_S_0_L_6_out : std_logic := '0'; 
signal C_78_S_0_L_7_out : std_logic := '0'; 
signal C_78_S_1_L_0_out : std_logic := '0'; 
signal C_78_S_1_L_1_out : std_logic := '0'; 
signal C_78_S_1_L_2_out : std_logic := '0'; 
signal C_78_S_1_L_3_out : std_logic := '0'; 
signal C_78_S_1_L_4_out : std_logic := '0'; 
signal C_78_S_1_L_5_out : std_logic := '0'; 
signal C_78_S_1_L_6_out : std_logic := '0'; 
signal C_78_S_1_L_7_out : std_logic := '0'; 
signal C_78_S_2_L_0_out : std_logic := '0'; 
signal C_78_S_2_L_1_out : std_logic := '0'; 
signal C_78_S_2_L_2_out : std_logic := '0'; 
signal C_78_S_2_L_3_out : std_logic := '0'; 
signal C_78_S_2_L_4_out : std_logic := '0'; 
signal C_78_S_2_L_5_out : std_logic := '0'; 
signal C_78_S_2_L_6_out : std_logic := '0'; 
signal C_78_S_2_L_7_out : std_logic := '0'; 
signal C_78_S_3_L_0_out : std_logic := '0'; 
signal C_78_S_3_L_1_out : std_logic := '0'; 
signal C_78_S_3_L_2_out : std_logic := '0'; 
signal C_78_S_3_L_3_out : std_logic := '0'; 
signal C_78_S_3_L_4_out : std_logic := '0'; 
signal C_78_S_3_L_5_out : std_logic := '0'; 
signal C_78_S_3_L_6_out : std_logic := '0'; 
signal C_78_S_3_L_7_out : std_logic := '0'; 
signal C_78_S_4_L_0_out : std_logic := '0'; 
signal C_78_S_4_L_1_out : std_logic := '0'; 
signal C_78_S_4_L_2_out : std_logic := '0'; 
signal C_78_S_4_L_3_out : std_logic := '0'; 
signal C_78_S_4_L_4_out : std_logic := '0'; 
signal C_78_S_4_L_5_out : std_logic := '0'; 
signal C_78_S_4_L_6_out : std_logic := '0'; 
signal C_78_S_4_L_7_out : std_logic := '0'; 
signal C_79_S_0_L_0_out : std_logic := '0'; 
signal C_79_S_0_L_1_out : std_logic := '0'; 
signal C_79_S_0_L_2_out : std_logic := '0'; 
signal C_79_S_0_L_3_out : std_logic := '0'; 
signal C_79_S_0_L_4_out : std_logic := '0'; 
signal C_79_S_0_L_5_out : std_logic := '0'; 
signal C_79_S_0_L_6_out : std_logic := '0'; 
signal C_79_S_0_L_7_out : std_logic := '0'; 
signal C_79_S_1_L_0_out : std_logic := '0'; 
signal C_79_S_1_L_1_out : std_logic := '0'; 
signal C_79_S_1_L_2_out : std_logic := '0'; 
signal C_79_S_1_L_3_out : std_logic := '0'; 
signal C_79_S_1_L_4_out : std_logic := '0'; 
signal C_79_S_1_L_5_out : std_logic := '0'; 
signal C_79_S_1_L_6_out : std_logic := '0'; 
signal C_79_S_1_L_7_out : std_logic := '0'; 
signal C_79_S_2_L_0_out : std_logic := '0'; 
signal C_79_S_2_L_1_out : std_logic := '0'; 
signal C_79_S_2_L_2_out : std_logic := '0'; 
signal C_79_S_2_L_3_out : std_logic := '0'; 
signal C_79_S_2_L_4_out : std_logic := '0'; 
signal C_79_S_2_L_5_out : std_logic := '0'; 
signal C_79_S_2_L_6_out : std_logic := '0'; 
signal C_79_S_2_L_7_out : std_logic := '0'; 
signal C_79_S_3_L_0_out : std_logic := '0'; 
signal C_79_S_3_L_1_out : std_logic := '0'; 
signal C_79_S_3_L_2_out : std_logic := '0'; 
signal C_79_S_3_L_3_out : std_logic := '0'; 
signal C_79_S_3_L_4_out : std_logic := '0'; 
signal C_79_S_3_L_5_out : std_logic := '0'; 
signal C_79_S_3_L_6_out : std_logic := '0'; 
signal C_79_S_3_L_7_out : std_logic := '0'; 
signal C_79_S_4_L_0_out : std_logic := '0'; 
signal C_79_S_4_L_1_out : std_logic := '0'; 
signal C_79_S_4_L_2_out : std_logic := '0'; 
signal C_79_S_4_L_3_out : std_logic := '0'; 
signal C_79_S_4_L_4_out : std_logic := '0'; 
signal C_79_S_4_L_5_out : std_logic := '0'; 
signal C_79_S_4_L_6_out : std_logic := '0'; 
signal C_79_S_4_L_7_out : std_logic := '0'; 

signal C_0_S_0_out : std_logic := '0'; 
signal C_0_S_1_out : std_logic := '0'; 
signal C_0_S_2_out : std_logic := '0'; 
signal C_0_S_3_out : std_logic := '0'; 
signal C_0_S_4_out : std_logic := '0'; 
signal C_1_S_0_out : std_logic := '0'; 
signal C_1_S_1_out : std_logic := '0'; 
signal C_1_S_2_out : std_logic := '0'; 
signal C_1_S_3_out : std_logic := '0'; 
signal C_1_S_4_out : std_logic := '0'; 
signal C_2_S_0_out : std_logic := '0'; 
signal C_2_S_1_out : std_logic := '0'; 
signal C_2_S_2_out : std_logic := '0'; 
signal C_2_S_3_out : std_logic := '0'; 
signal C_2_S_4_out : std_logic := '0'; 
signal C_3_S_0_out : std_logic := '0'; 
signal C_3_S_1_out : std_logic := '0'; 
signal C_3_S_2_out : std_logic := '0'; 
signal C_3_S_3_out : std_logic := '0'; 
signal C_3_S_4_out : std_logic := '0'; 
signal C_4_S_0_out : std_logic := '0'; 
signal C_4_S_1_out : std_logic := '0'; 
signal C_4_S_2_out : std_logic := '0'; 
signal C_4_S_3_out : std_logic := '0'; 
signal C_4_S_4_out : std_logic := '0'; 
signal C_5_S_0_out : std_logic := '0'; 
signal C_5_S_1_out : std_logic := '0'; 
signal C_5_S_2_out : std_logic := '0'; 
signal C_5_S_3_out : std_logic := '0'; 
signal C_5_S_4_out : std_logic := '0'; 
signal C_6_S_0_out : std_logic := '0'; 
signal C_6_S_1_out : std_logic := '0'; 
signal C_6_S_2_out : std_logic := '0'; 
signal C_6_S_3_out : std_logic := '0'; 
signal C_6_S_4_out : std_logic := '0'; 
signal C_7_S_0_out : std_logic := '0'; 
signal C_7_S_1_out : std_logic := '0'; 
signal C_7_S_2_out : std_logic := '0'; 
signal C_7_S_3_out : std_logic := '0'; 
signal C_7_S_4_out : std_logic := '0'; 
signal C_8_S_0_out : std_logic := '0'; 
signal C_8_S_1_out : std_logic := '0'; 
signal C_8_S_2_out : std_logic := '0'; 
signal C_8_S_3_out : std_logic := '0'; 
signal C_8_S_4_out : std_logic := '0'; 
signal C_9_S_0_out : std_logic := '0'; 
signal C_9_S_1_out : std_logic := '0'; 
signal C_9_S_2_out : std_logic := '0'; 
signal C_9_S_3_out : std_logic := '0'; 
signal C_9_S_4_out : std_logic := '0'; 
signal C_10_S_0_out : std_logic := '0'; 
signal C_10_S_1_out : std_logic := '0'; 
signal C_10_S_2_out : std_logic := '0'; 
signal C_10_S_3_out : std_logic := '0'; 
signal C_10_S_4_out : std_logic := '0'; 
signal C_11_S_0_out : std_logic := '0'; 
signal C_11_S_1_out : std_logic := '0'; 
signal C_11_S_2_out : std_logic := '0'; 
signal C_11_S_3_out : std_logic := '0'; 
signal C_11_S_4_out : std_logic := '0'; 
signal C_12_S_0_out : std_logic := '0'; 
signal C_12_S_1_out : std_logic := '0'; 
signal C_12_S_2_out : std_logic := '0'; 
signal C_12_S_3_out : std_logic := '0'; 
signal C_12_S_4_out : std_logic := '0'; 
signal C_13_S_0_out : std_logic := '0'; 
signal C_13_S_1_out : std_logic := '0'; 
signal C_13_S_2_out : std_logic := '0'; 
signal C_13_S_3_out : std_logic := '0'; 
signal C_13_S_4_out : std_logic := '0'; 
signal C_14_S_0_out : std_logic := '0'; 
signal C_14_S_1_out : std_logic := '0'; 
signal C_14_S_2_out : std_logic := '0'; 
signal C_14_S_3_out : std_logic := '0'; 
signal C_14_S_4_out : std_logic := '0'; 
signal C_15_S_0_out : std_logic := '0'; 
signal C_15_S_1_out : std_logic := '0'; 
signal C_15_S_2_out : std_logic := '0'; 
signal C_15_S_3_out : std_logic := '0'; 
signal C_15_S_4_out : std_logic := '0'; 
signal C_16_S_0_out : std_logic := '0'; 
signal C_16_S_1_out : std_logic := '0'; 
signal C_16_S_2_out : std_logic := '0'; 
signal C_16_S_3_out : std_logic := '0'; 
signal C_16_S_4_out : std_logic := '0'; 
signal C_17_S_0_out : std_logic := '0'; 
signal C_17_S_1_out : std_logic := '0'; 
signal C_17_S_2_out : std_logic := '0'; 
signal C_17_S_3_out : std_logic := '0'; 
signal C_17_S_4_out : std_logic := '0'; 
signal C_18_S_0_out : std_logic := '0'; 
signal C_18_S_1_out : std_logic := '0'; 
signal C_18_S_2_out : std_logic := '0'; 
signal C_18_S_3_out : std_logic := '0'; 
signal C_18_S_4_out : std_logic := '0'; 
signal C_19_S_0_out : std_logic := '0'; 
signal C_19_S_1_out : std_logic := '0'; 
signal C_19_S_2_out : std_logic := '0'; 
signal C_19_S_3_out : std_logic := '0'; 
signal C_19_S_4_out : std_logic := '0'; 
signal C_20_S_0_out : std_logic := '0'; 
signal C_20_S_1_out : std_logic := '0'; 
signal C_20_S_2_out : std_logic := '0'; 
signal C_20_S_3_out : std_logic := '0'; 
signal C_20_S_4_out : std_logic := '0'; 
signal C_21_S_0_out : std_logic := '0'; 
signal C_21_S_1_out : std_logic := '0'; 
signal C_21_S_2_out : std_logic := '0'; 
signal C_21_S_3_out : std_logic := '0'; 
signal C_21_S_4_out : std_logic := '0'; 
signal C_22_S_0_out : std_logic := '0'; 
signal C_22_S_1_out : std_logic := '0'; 
signal C_22_S_2_out : std_logic := '0'; 
signal C_22_S_3_out : std_logic := '0'; 
signal C_22_S_4_out : std_logic := '0'; 
signal C_23_S_0_out : std_logic := '0'; 
signal C_23_S_1_out : std_logic := '0'; 
signal C_23_S_2_out : std_logic := '0'; 
signal C_23_S_3_out : std_logic := '0'; 
signal C_23_S_4_out : std_logic := '0'; 
signal C_24_S_0_out : std_logic := '0'; 
signal C_24_S_1_out : std_logic := '0'; 
signal C_24_S_2_out : std_logic := '0'; 
signal C_24_S_3_out : std_logic := '0'; 
signal C_24_S_4_out : std_logic := '0'; 
signal C_25_S_0_out : std_logic := '0'; 
signal C_25_S_1_out : std_logic := '0'; 
signal C_25_S_2_out : std_logic := '0'; 
signal C_25_S_3_out : std_logic := '0'; 
signal C_25_S_4_out : std_logic := '0'; 
signal C_26_S_0_out : std_logic := '0'; 
signal C_26_S_1_out : std_logic := '0'; 
signal C_26_S_2_out : std_logic := '0'; 
signal C_26_S_3_out : std_logic := '0'; 
signal C_26_S_4_out : std_logic := '0'; 
signal C_27_S_0_out : std_logic := '0'; 
signal C_27_S_1_out : std_logic := '0'; 
signal C_27_S_2_out : std_logic := '0'; 
signal C_27_S_3_out : std_logic := '0'; 
signal C_27_S_4_out : std_logic := '0'; 
signal C_28_S_0_out : std_logic := '0'; 
signal C_28_S_1_out : std_logic := '0'; 
signal C_28_S_2_out : std_logic := '0'; 
signal C_28_S_3_out : std_logic := '0'; 
signal C_28_S_4_out : std_logic := '0'; 
signal C_29_S_0_out : std_logic := '0'; 
signal C_29_S_1_out : std_logic := '0'; 
signal C_29_S_2_out : std_logic := '0'; 
signal C_29_S_3_out : std_logic := '0'; 
signal C_29_S_4_out : std_logic := '0'; 
signal C_30_S_0_out : std_logic := '0'; 
signal C_30_S_1_out : std_logic := '0'; 
signal C_30_S_2_out : std_logic := '0'; 
signal C_30_S_3_out : std_logic := '0'; 
signal C_30_S_4_out : std_logic := '0'; 
signal C_31_S_0_out : std_logic := '0'; 
signal C_31_S_1_out : std_logic := '0'; 
signal C_31_S_2_out : std_logic := '0'; 
signal C_31_S_3_out : std_logic := '0'; 
signal C_31_S_4_out : std_logic := '0'; 
signal C_32_S_0_out : std_logic := '0'; 
signal C_32_S_1_out : std_logic := '0'; 
signal C_32_S_2_out : std_logic := '0'; 
signal C_32_S_3_out : std_logic := '0'; 
signal C_32_S_4_out : std_logic := '0'; 
signal C_33_S_0_out : std_logic := '0'; 
signal C_33_S_1_out : std_logic := '0'; 
signal C_33_S_2_out : std_logic := '0'; 
signal C_33_S_3_out : std_logic := '0'; 
signal C_33_S_4_out : std_logic := '0'; 
signal C_34_S_0_out : std_logic := '0'; 
signal C_34_S_1_out : std_logic := '0'; 
signal C_34_S_2_out : std_logic := '0'; 
signal C_34_S_3_out : std_logic := '0'; 
signal C_34_S_4_out : std_logic := '0'; 
signal C_35_S_0_out : std_logic := '0'; 
signal C_35_S_1_out : std_logic := '0'; 
signal C_35_S_2_out : std_logic := '0'; 
signal C_35_S_3_out : std_logic := '0'; 
signal C_35_S_4_out : std_logic := '0'; 
signal C_36_S_0_out : std_logic := '0'; 
signal C_36_S_1_out : std_logic := '0'; 
signal C_36_S_2_out : std_logic := '0'; 
signal C_36_S_3_out : std_logic := '0'; 
signal C_36_S_4_out : std_logic := '0'; 
signal C_37_S_0_out : std_logic := '0'; 
signal C_37_S_1_out : std_logic := '0'; 
signal C_37_S_2_out : std_logic := '0'; 
signal C_37_S_3_out : std_logic := '0'; 
signal C_37_S_4_out : std_logic := '0'; 
signal C_38_S_0_out : std_logic := '0'; 
signal C_38_S_1_out : std_logic := '0'; 
signal C_38_S_2_out : std_logic := '0'; 
signal C_38_S_3_out : std_logic := '0'; 
signal C_38_S_4_out : std_logic := '0'; 
signal C_39_S_0_out : std_logic := '0'; 
signal C_39_S_1_out : std_logic := '0'; 
signal C_39_S_2_out : std_logic := '0'; 
signal C_39_S_3_out : std_logic := '0'; 
signal C_39_S_4_out : std_logic := '0'; 
signal C_40_S_0_out : std_logic := '0'; 
signal C_40_S_1_out : std_logic := '0'; 
signal C_40_S_2_out : std_logic := '0'; 
signal C_40_S_3_out : std_logic := '0'; 
signal C_40_S_4_out : std_logic := '0'; 
signal C_41_S_0_out : std_logic := '0'; 
signal C_41_S_1_out : std_logic := '0'; 
signal C_41_S_2_out : std_logic := '0'; 
signal C_41_S_3_out : std_logic := '0'; 
signal C_41_S_4_out : std_logic := '0'; 
signal C_42_S_0_out : std_logic := '0'; 
signal C_42_S_1_out : std_logic := '0'; 
signal C_42_S_2_out : std_logic := '0'; 
signal C_42_S_3_out : std_logic := '0'; 
signal C_42_S_4_out : std_logic := '0'; 
signal C_43_S_0_out : std_logic := '0'; 
signal C_43_S_1_out : std_logic := '0'; 
signal C_43_S_2_out : std_logic := '0'; 
signal C_43_S_3_out : std_logic := '0'; 
signal C_43_S_4_out : std_logic := '0'; 
signal C_44_S_0_out : std_logic := '0'; 
signal C_44_S_1_out : std_logic := '0'; 
signal C_44_S_2_out : std_logic := '0'; 
signal C_44_S_3_out : std_logic := '0'; 
signal C_44_S_4_out : std_logic := '0'; 
signal C_45_S_0_out : std_logic := '0'; 
signal C_45_S_1_out : std_logic := '0'; 
signal C_45_S_2_out : std_logic := '0'; 
signal C_45_S_3_out : std_logic := '0'; 
signal C_45_S_4_out : std_logic := '0'; 
signal C_46_S_0_out : std_logic := '0'; 
signal C_46_S_1_out : std_logic := '0'; 
signal C_46_S_2_out : std_logic := '0'; 
signal C_46_S_3_out : std_logic := '0'; 
signal C_46_S_4_out : std_logic := '0'; 
signal C_47_S_0_out : std_logic := '0'; 
signal C_47_S_1_out : std_logic := '0'; 
signal C_47_S_2_out : std_logic := '0'; 
signal C_47_S_3_out : std_logic := '0'; 
signal C_47_S_4_out : std_logic := '0'; 
signal C_48_S_0_out : std_logic := '0'; 
signal C_48_S_1_out : std_logic := '0'; 
signal C_48_S_2_out : std_logic := '0'; 
signal C_48_S_3_out : std_logic := '0'; 
signal C_48_S_4_out : std_logic := '0'; 
signal C_49_S_0_out : std_logic := '0'; 
signal C_49_S_1_out : std_logic := '0'; 
signal C_49_S_2_out : std_logic := '0'; 
signal C_49_S_3_out : std_logic := '0'; 
signal C_49_S_4_out : std_logic := '0'; 
signal C_50_S_0_out : std_logic := '0'; 
signal C_50_S_1_out : std_logic := '0'; 
signal C_50_S_2_out : std_logic := '0'; 
signal C_50_S_3_out : std_logic := '0'; 
signal C_50_S_4_out : std_logic := '0'; 
signal C_51_S_0_out : std_logic := '0'; 
signal C_51_S_1_out : std_logic := '0'; 
signal C_51_S_2_out : std_logic := '0'; 
signal C_51_S_3_out : std_logic := '0'; 
signal C_51_S_4_out : std_logic := '0'; 
signal C_52_S_0_out : std_logic := '0'; 
signal C_52_S_1_out : std_logic := '0'; 
signal C_52_S_2_out : std_logic := '0'; 
signal C_52_S_3_out : std_logic := '0'; 
signal C_52_S_4_out : std_logic := '0'; 
signal C_53_S_0_out : std_logic := '0'; 
signal C_53_S_1_out : std_logic := '0'; 
signal C_53_S_2_out : std_logic := '0'; 
signal C_53_S_3_out : std_logic := '0'; 
signal C_53_S_4_out : std_logic := '0'; 
signal C_54_S_0_out : std_logic := '0'; 
signal C_54_S_1_out : std_logic := '0'; 
signal C_54_S_2_out : std_logic := '0'; 
signal C_54_S_3_out : std_logic := '0'; 
signal C_54_S_4_out : std_logic := '0'; 
signal C_55_S_0_out : std_logic := '0'; 
signal C_55_S_1_out : std_logic := '0'; 
signal C_55_S_2_out : std_logic := '0'; 
signal C_55_S_3_out : std_logic := '0'; 
signal C_55_S_4_out : std_logic := '0'; 
signal C_56_S_0_out : std_logic := '0'; 
signal C_56_S_1_out : std_logic := '0'; 
signal C_56_S_2_out : std_logic := '0'; 
signal C_56_S_3_out : std_logic := '0'; 
signal C_56_S_4_out : std_logic := '0'; 
signal C_57_S_0_out : std_logic := '0'; 
signal C_57_S_1_out : std_logic := '0'; 
signal C_57_S_2_out : std_logic := '0'; 
signal C_57_S_3_out : std_logic := '0'; 
signal C_57_S_4_out : std_logic := '0'; 
signal C_58_S_0_out : std_logic := '0'; 
signal C_58_S_1_out : std_logic := '0'; 
signal C_58_S_2_out : std_logic := '0'; 
signal C_58_S_3_out : std_logic := '0'; 
signal C_58_S_4_out : std_logic := '0'; 
signal C_59_S_0_out : std_logic := '0'; 
signal C_59_S_1_out : std_logic := '0'; 
signal C_59_S_2_out : std_logic := '0'; 
signal C_59_S_3_out : std_logic := '0'; 
signal C_59_S_4_out : std_logic := '0'; 
signal C_60_S_0_out : std_logic := '0'; 
signal C_60_S_1_out : std_logic := '0'; 
signal C_60_S_2_out : std_logic := '0'; 
signal C_60_S_3_out : std_logic := '0'; 
signal C_60_S_4_out : std_logic := '0'; 
signal C_61_S_0_out : std_logic := '0'; 
signal C_61_S_1_out : std_logic := '0'; 
signal C_61_S_2_out : std_logic := '0'; 
signal C_61_S_3_out : std_logic := '0'; 
signal C_61_S_4_out : std_logic := '0'; 
signal C_62_S_0_out : std_logic := '0'; 
signal C_62_S_1_out : std_logic := '0'; 
signal C_62_S_2_out : std_logic := '0'; 
signal C_62_S_3_out : std_logic := '0'; 
signal C_62_S_4_out : std_logic := '0'; 
signal C_63_S_0_out : std_logic := '0'; 
signal C_63_S_1_out : std_logic := '0'; 
signal C_63_S_2_out : std_logic := '0'; 
signal C_63_S_3_out : std_logic := '0'; 
signal C_63_S_4_out : std_logic := '0'; 
signal C_64_S_0_out : std_logic := '0'; 
signal C_64_S_1_out : std_logic := '0'; 
signal C_64_S_2_out : std_logic := '0'; 
signal C_64_S_3_out : std_logic := '0'; 
signal C_64_S_4_out : std_logic := '0'; 
signal C_65_S_0_out : std_logic := '0'; 
signal C_65_S_1_out : std_logic := '0'; 
signal C_65_S_2_out : std_logic := '0'; 
signal C_65_S_3_out : std_logic := '0'; 
signal C_65_S_4_out : std_logic := '0'; 
signal C_66_S_0_out : std_logic := '0'; 
signal C_66_S_1_out : std_logic := '0'; 
signal C_66_S_2_out : std_logic := '0'; 
signal C_66_S_3_out : std_logic := '0'; 
signal C_66_S_4_out : std_logic := '0'; 
signal C_67_S_0_out : std_logic := '0'; 
signal C_67_S_1_out : std_logic := '0'; 
signal C_67_S_2_out : std_logic := '0'; 
signal C_67_S_3_out : std_logic := '0'; 
signal C_67_S_4_out : std_logic := '0'; 
signal C_68_S_0_out : std_logic := '0'; 
signal C_68_S_1_out : std_logic := '0'; 
signal C_68_S_2_out : std_logic := '0'; 
signal C_68_S_3_out : std_logic := '0'; 
signal C_68_S_4_out : std_logic := '0'; 
signal C_69_S_0_out : std_logic := '0'; 
signal C_69_S_1_out : std_logic := '0'; 
signal C_69_S_2_out : std_logic := '0'; 
signal C_69_S_3_out : std_logic := '0'; 
signal C_69_S_4_out : std_logic := '0'; 
signal C_70_S_0_out : std_logic := '0'; 
signal C_70_S_1_out : std_logic := '0'; 
signal C_70_S_2_out : std_logic := '0'; 
signal C_70_S_3_out : std_logic := '0'; 
signal C_70_S_4_out : std_logic := '0'; 
signal C_71_S_0_out : std_logic := '0'; 
signal C_71_S_1_out : std_logic := '0'; 
signal C_71_S_2_out : std_logic := '0'; 
signal C_71_S_3_out : std_logic := '0'; 
signal C_71_S_4_out : std_logic := '0'; 
signal C_72_S_0_out : std_logic := '0'; 
signal C_72_S_1_out : std_logic := '0'; 
signal C_72_S_2_out : std_logic := '0'; 
signal C_72_S_3_out : std_logic := '0'; 
signal C_72_S_4_out : std_logic := '0'; 
signal C_73_S_0_out : std_logic := '0'; 
signal C_73_S_1_out : std_logic := '0'; 
signal C_73_S_2_out : std_logic := '0'; 
signal C_73_S_3_out : std_logic := '0'; 
signal C_73_S_4_out : std_logic := '0'; 
signal C_74_S_0_out : std_logic := '0'; 
signal C_74_S_1_out : std_logic := '0'; 
signal C_74_S_2_out : std_logic := '0'; 
signal C_74_S_3_out : std_logic := '0'; 
signal C_74_S_4_out : std_logic := '0'; 
signal C_75_S_0_out : std_logic := '0'; 
signal C_75_S_1_out : std_logic := '0'; 
signal C_75_S_2_out : std_logic := '0'; 
signal C_75_S_3_out : std_logic := '0'; 
signal C_75_S_4_out : std_logic := '0'; 
signal C_76_S_0_out : std_logic := '0'; 
signal C_76_S_1_out : std_logic := '0'; 
signal C_76_S_2_out : std_logic := '0'; 
signal C_76_S_3_out : std_logic := '0'; 
signal C_76_S_4_out : std_logic := '0'; 
signal C_77_S_0_out : std_logic := '0'; 
signal C_77_S_1_out : std_logic := '0'; 
signal C_77_S_2_out : std_logic := '0'; 
signal C_77_S_3_out : std_logic := '0'; 
signal C_77_S_4_out : std_logic := '0'; 
signal C_78_S_0_out : std_logic := '0'; 
signal C_78_S_1_out : std_logic := '0'; 
signal C_78_S_2_out : std_logic := '0'; 
signal C_78_S_3_out : std_logic := '0'; 
signal C_78_S_4_out : std_logic := '0'; 
signal C_79_S_0_out : std_logic := '0'; 
signal C_79_S_1_out : std_logic := '0'; 
signal C_79_S_2_out : std_logic := '0'; 
signal C_79_S_3_out : std_logic := '0'; 
signal C_79_S_4_out : std_logic := '0'; 
begin

C_0_S_0_L_0_inst : LUT8 generic map(INIT => "1111111011101110101011100000000001110000000000001010000000110000000011000100000010101010010000000000000000000000000000000000000011101110000001001010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_0_L_0_out, I0 =>  inp_feat(446), I1 =>  inp_feat(110), I2 =>  inp_feat(509), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_0_S_0_L_1_inst : LUT8 generic map(INIT => "0111000110100010101001001010000000010101000000001010010000000000111111111010101010111111000000000010000000000010100011000000000010110101101000001011010111110000000101110000000000011111000000001001000100000000101101011010000000010101000000000000010100000000") port map( O =>C_0_S_0_L_1_out, I0 =>  inp_feat(348), I1 =>  inp_feat(323), I2 =>  inp_feat(508), I3 =>  inp_feat(72), I4 =>  inp_feat(329), I5 =>  inp_feat(282), I6 =>  inp_feat(293), I7 =>  inp_feat(15)); 
C_0_S_0_L_2_inst : LUT8 generic map(INIT => "0010001011100010111010101010101011100000111000001000000011000000101000001110000010100000100000001100000011000000100000001100000000100000000000000010000000100000100000001100000010000000110000001010000010000000101000001000000010000000110000001100000011000000") port map( O =>C_0_S_0_L_2_out, I0 =>  inp_feat(282), I1 =>  inp_feat(72), I2 =>  inp_feat(22), I3 =>  inp_feat(302), I4 =>  inp_feat(41), I5 =>  inp_feat(9), I6 =>  inp_feat(71), I7 =>  inp_feat(152)); 
C_0_S_0_L_3_inst : LUT8 generic map(INIT => "1110110010101100011011100000111000010001000000100000100000000000111111001111010100001100000011010110110100000111001011100000111010001000100010100000001100001000001011100000000000000000000000001000101000000100000010100000100011111111000010110010101000000010") port map( O =>C_0_S_0_L_3_out, I0 =>  inp_feat(483), I1 =>  inp_feat(100), I2 =>  inp_feat(323), I3 =>  inp_feat(238), I4 =>  inp_feat(49), I5 =>  inp_feat(462), I6 =>  inp_feat(478), I7 =>  inp_feat(15)); 
C_0_S_0_L_4_inst : LUT8 generic map(INIT => "0010111010101000000000011000000010100000101000000000000000100000111111111011101000011001000000000010000010000000000000000000000011101110101110101111000110110001001010101010101010000000101000001111101011111010101100010111000010100010101010100000000000000000") port map( O =>C_0_S_0_L_4_out, I0 =>  inp_feat(170), I1 =>  inp_feat(11), I2 =>  inp_feat(499), I3 =>  inp_feat(317), I4 =>  inp_feat(269), I5 =>  inp_feat(149), I6 =>  inp_feat(323), I7 =>  inp_feat(478)); 
C_0_S_0_L_5_inst : LUT8 generic map(INIT => "0111000111110111101010000000000000000000000000001000100000000000111100111111011010101010000000000000000000000000100000000000000011110000000000001111100000000000000000000000000010001000000000001110000000000000111100000000000000000000000000001000000000000000") port map( O =>C_0_S_0_L_5_out, I0 =>  inp_feat(10), I1 =>  inp_feat(71), I2 =>  inp_feat(390), I3 =>  inp_feat(281), I4 =>  inp_feat(415), I5 =>  inp_feat(122), I6 =>  inp_feat(108), I7 =>  inp_feat(235)); 
C_0_S_0_L_6_inst : LUT8 generic map(INIT => "0100110000001000110010100000000011111100000000001100101000001000110011000000000010000000000000001111100000000000000000000000000011101100000010001000100000000000110010000000000000001000000000001000000000000000101000000000000000100000000000000000000000000000") port map( O =>C_0_S_0_L_6_out, I0 =>  inp_feat(222), I1 =>  inp_feat(463), I2 =>  inp_feat(128), I3 =>  inp_feat(498), I4 =>  inp_feat(198), I5 =>  inp_feat(372), I6 =>  inp_feat(360), I7 =>  inp_feat(58)); 
C_0_S_0_L_7_inst : LUT8 generic map(INIT => "0010111111111111111111001100010011011101110011000000000000000000101010001111010010000000010001001000000000000000000000000000000010111111001011111011101000000000101100110000110000000000000000000010000010100000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_0_L_7_out, I0 =>  inp_feat(195), I1 =>  inp_feat(293), I2 =>  inp_feat(15), I3 =>  inp_feat(496), I4 =>  inp_feat(360), I5 =>  inp_feat(304), I6 =>  inp_feat(446), I7 =>  inp_feat(288)); 
C_0_S_1_L_0_inst : LUT8 generic map(INIT => "1111111011101110101011100000000001110000000000001010000000110000000011000100000010101010010000000000000000000000000000000000000011101110000001001010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_1_L_0_out, I0 =>  inp_feat(446), I1 =>  inp_feat(110), I2 =>  inp_feat(509), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_0_S_1_L_1_inst : LUT8 generic map(INIT => "0010010011110010111101011101000001100001000000001111000100000000111111011110101001000101000000000010000000000010010001010000000011110101110100001101010111010000011101010000000001010001000000000100010100000000010001010100000001110101000000000000010100000000") port map( O =>C_0_S_1_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(289), I2 =>  inp_feat(508), I3 =>  inp_feat(72), I4 =>  inp_feat(329), I5 =>  inp_feat(282), I6 =>  inp_feat(293), I7 =>  inp_feat(15)); 
C_0_S_1_L_2_inst : LUT8 generic map(INIT => "0001001011100010111010001111000010101010101000101100100010000000100000000100000011001000000000001100000000000000110000000000000011111000100001011010100001011101100010001000000000001000000000011100100011000000100000000000000010000000100000000000000000000000") port map( O =>C_0_S_1_L_2_out, I0 =>  inp_feat(338), I1 =>  inp_feat(11), I2 =>  inp_feat(82), I3 =>  inp_feat(354), I4 =>  inp_feat(243), I5 =>  inp_feat(500), I6 =>  inp_feat(360), I7 =>  inp_feat(478)); 
C_0_S_1_L_3_inst : LUT8 generic map(INIT => "1101000010000000000000001000000010001000100010000000000010000000111100001000000010000000100000001110100010001000100000001000100010101010101000101110000010100000100010000000000000000000000000001111000000000000100000001000000011101000000000001000000010000000") port map( O =>C_0_S_1_L_3_out, I0 =>  inp_feat(276), I1 =>  inp_feat(260), I2 =>  inp_feat(359), I3 =>  inp_feat(353), I4 =>  inp_feat(440), I5 =>  inp_feat(64), I6 =>  inp_feat(15), I7 =>  inp_feat(71)); 
C_0_S_1_L_4_inst : LUT8 generic map(INIT => "0100000011100111111100101010111111111100101011111111100011101110110000001100000010100000100000001010000000000000101000000000000010000000000000001010000010000000000000000000000010100000000000000000000010000000100000001000000000000000000000000000000000000000") port map( O =>C_0_S_1_L_4_out, I0 =>  inp_feat(280), I1 =>  inp_feat(295), I2 =>  inp_feat(282), I3 =>  inp_feat(302), I4 =>  inp_feat(71), I5 =>  inp_feat(351), I6 =>  inp_feat(72), I7 =>  inp_feat(147)); 
C_0_S_1_L_5_inst : LUT8 generic map(INIT => "1011001011110100111100101111000000000000110000001111100111110000001001101110000000100000000000000000000000000000000000000000000011110010111101000011101001010000000000000100000000010000010100001111011111110111000000000000000000000000000000000000000000000000") port map( O =>C_0_S_1_L_5_out, I0 =>  inp_feat(172), I1 =>  inp_feat(365), I2 =>  inp_feat(260), I3 =>  inp_feat(154), I4 =>  inp_feat(90), I5 =>  inp_feat(369), I6 =>  inp_feat(312), I7 =>  inp_feat(323)); 
C_0_S_1_L_6_inst : LUT8 generic map(INIT => "0010111010001000111011100010101011101000110010001100100010101010000000000000000000000000000000001010000000000000000000000000000011111010100010001100100010001000111010001100100011101000100010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_1_L_6_out, I0 =>  inp_feat(164), I1 =>  inp_feat(238), I2 =>  inp_feat(301), I3 =>  inp_feat(378), I4 =>  inp_feat(195), I5 =>  inp_feat(293), I6 =>  inp_feat(70), I7 =>  inp_feat(41)); 
C_0_S_1_L_7_inst : LUT8 generic map(INIT => "1010101011111010101010001010000000001000001000001010100000100000001000000000000000001000000000000000100000000000000010000000000000101010101011100000001000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_1_L_7_out, I0 =>  inp_feat(70), I1 =>  inp_feat(297), I2 =>  inp_feat(86), I3 =>  inp_feat(293), I4 =>  inp_feat(446), I5 =>  inp_feat(258), I6 =>  inp_feat(122), I7 =>  inp_feat(338)); 
C_0_S_2_L_0_inst : LUT8 generic map(INIT => "1111111011101110101011100000000001110000000000001010000000110000000011000100000010101010010000000000000000000000000000000000000011101110000001001010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_2_L_0_out, I0 =>  inp_feat(446), I1 =>  inp_feat(110), I2 =>  inp_feat(509), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_0_S_2_L_1_inst : LUT8 generic map(INIT => "0010010011110010111101011101000001100001000000001111000100000000111111011110101001000101000000000010000000000010010001010000000011110101110100001101010111010000011101010000000001010001000000000100010100000000010001010100000001110101000000000000010100000000") port map( O =>C_0_S_2_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(289), I2 =>  inp_feat(508), I3 =>  inp_feat(72), I4 =>  inp_feat(329), I5 =>  inp_feat(282), I6 =>  inp_feat(293), I7 =>  inp_feat(15)); 
C_0_S_2_L_2_inst : LUT8 generic map(INIT => "0001001011100010111010001111000010101010101000101100100010000000100000000100000011001000000000001100000000000000110000000000000011111000100001011010100001011101100010001000000000001000000000011100100011000000100000000000000010000000100000000000000000000000") port map( O =>C_0_S_2_L_2_out, I0 =>  inp_feat(338), I1 =>  inp_feat(11), I2 =>  inp_feat(82), I3 =>  inp_feat(354), I4 =>  inp_feat(243), I5 =>  inp_feat(500), I6 =>  inp_feat(360), I7 =>  inp_feat(478)); 
C_0_S_2_L_3_inst : LUT8 generic map(INIT => "1001101011001000000010000000000010100010100000000000000010100000111000001100000010000000100000001010101010000000101010001000000010100010101000001000100010001000100000000000000000000000000000001010000010000000100000000010000010100010000000001000000000000000") port map( O =>C_0_S_2_L_3_out, I0 =>  inp_feat(150), I1 =>  inp_feat(7), I2 =>  inp_feat(446), I3 =>  inp_feat(238), I4 =>  inp_feat(440), I5 =>  inp_feat(64), I6 =>  inp_feat(15), I7 =>  inp_feat(71)); 
C_0_S_2_L_4_inst : LUT8 generic map(INIT => "0110010011001000101010101010000011111101110111001011000110100000110011001100100010000000100000001101110111001100100000001000000011000000000010001000100010001000101000010000000000000000000000001000000010000000001000000000000010100000110000000000000000000000") port map( O =>C_0_S_2_L_4_out, I0 =>  inp_feat(409), I1 =>  inp_feat(97), I2 =>  inp_feat(440), I3 =>  inp_feat(290), I4 =>  inp_feat(496), I5 =>  inp_feat(221), I6 =>  inp_feat(71), I7 =>  inp_feat(117)); 
C_0_S_2_L_5_inst : LUT8 generic map(INIT => "1110110111001111110010000010000000000000000000000000100000000000110011101010111011001000101010001000000000001000000010000000100000101000000000000100000000000000000000000000000011001000000000001100000010000000110010001000100000000000100000001000100010000000") port map( O =>C_0_S_2_L_5_out, I0 =>  inp_feat(485), I1 =>  inp_feat(475), I2 =>  inp_feat(71), I3 =>  inp_feat(413), I4 =>  inp_feat(129), I5 =>  inp_feat(508), I6 =>  inp_feat(323), I7 =>  inp_feat(113)); 
C_0_S_2_L_6_inst : LUT8 generic map(INIT => "1000111011101110111010001000100000001100110011011000100010001000000000000000010010000000000000000000110000001100000000000000000011001110010000101100000010000000000000000000000010000000000000001100110000000000100000000000000000000000000000000000000000000000") port map( O =>C_0_S_2_L_6_out, I0 =>  inp_feat(130), I1 =>  inp_feat(193), I2 =>  inp_feat(302), I3 =>  inp_feat(451), I4 =>  inp_feat(293), I5 =>  inp_feat(508), I6 =>  inp_feat(85), I7 =>  inp_feat(229)); 
C_0_S_2_L_7_inst : LUT8 generic map(INIT => "0100110111001100000000000000000010100100110011000000000001000000110011001100010000000100000000000000000000000000000000000000000011111111110000000000000000000000110000001000000000000000000000001100100010000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_2_L_7_out, I0 =>  inp_feat(293), I1 =>  inp_feat(258), I2 =>  inp_feat(350), I3 =>  inp_feat(71), I4 =>  inp_feat(70), I5 =>  inp_feat(310), I6 =>  inp_feat(252), I7 =>  inp_feat(212)); 
C_0_S_3_L_0_inst : LUT8 generic map(INIT => "1111111011101110101011100000000001110000000000001010000000110000000011000100000010101010010000000000000000000000000000000000000011101110000001001010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_3_L_0_out, I0 =>  inp_feat(446), I1 =>  inp_feat(110), I2 =>  inp_feat(509), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_0_S_3_L_1_inst : LUT8 generic map(INIT => "0010010011110010111101011101000001100001000000001111000100000000111111011110101001000101000000000010000000000010010001010000000011110101110100001101010111010000011101010000000001010001000000000100010100000000010001010100000001110101000000000000010100000000") port map( O =>C_0_S_3_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(289), I2 =>  inp_feat(508), I3 =>  inp_feat(72), I4 =>  inp_feat(329), I5 =>  inp_feat(282), I6 =>  inp_feat(293), I7 =>  inp_feat(15)); 
C_0_S_3_L_2_inst : LUT8 generic map(INIT => "0100010100000000110010001000100011000101000000001111000010100000100000000000000001000000000000001100001000000000000000000000000011011011100000000000001110000100010100010000000000011111101010111101100110000000010000001000000010000000000000000000000000000000") port map( O =>C_0_S_3_L_2_out, I0 =>  inp_feat(391), I1 =>  inp_feat(378), I2 =>  inp_feat(82), I3 =>  inp_feat(234), I4 =>  inp_feat(354), I5 =>  inp_feat(243), I6 =>  inp_feat(360), I7 =>  inp_feat(478)); 
C_0_S_3_L_3_inst : LUT8 generic map(INIT => "0010111010110010111000101000001010101111101010001010100010000000110011000000000011001100000000000010000000000000000000000000000010100010101000001111001100000000010001110000000010010001000000000100000000000000110000000000000000000000000000000000000000000000") port map( O =>C_0_S_3_L_3_out, I0 =>  inp_feat(287), I1 =>  inp_feat(72), I2 =>  inp_feat(64), I3 =>  inp_feat(276), I4 =>  inp_feat(71), I5 =>  inp_feat(415), I6 =>  inp_feat(348), I7 =>  inp_feat(290)); 
C_0_S_3_L_4_inst : LUT8 generic map(INIT => "1110110100001101111111100100010101101100000000011111100000000101101010000000100011111011001110111000100010001000111010001000100000000000000010001010000000000000000000000000000000000000000000001000100000011000101110101010101100000000000000000000000000000000") port map( O =>C_0_S_3_L_4_out, I0 =>  inp_feat(436), I1 =>  inp_feat(505), I2 =>  inp_feat(272), I3 =>  inp_feat(390), I4 =>  inp_feat(478), I5 =>  inp_feat(435), I6 =>  inp_feat(302), I7 =>  inp_feat(282)); 
C_0_S_3_L_5_inst : LUT8 generic map(INIT => "1111111111111010001010101010001001010101111100000000000000000000100011111011101000000000001000000101010101111010000000000010000001001011011100100010000100100000010000010100000000010000000000000000000000000000000000000010000000000000000000000000000000000000") port map( O =>C_0_S_3_L_5_out, I0 =>  inp_feat(371), I1 =>  inp_feat(71), I2 =>  inp_feat(81), I3 =>  inp_feat(376), I4 =>  inp_feat(260), I5 =>  inp_feat(390), I6 =>  inp_feat(80), I7 =>  inp_feat(275)); 
C_0_S_3_L_6_inst : LUT8 generic map(INIT => "1100101001001111101010000000110111101010000010001101111000001100001000000000000010101000000000001010101000000000101010100000000000000000000000000000001000000000001010100000000000001010000000000010001000000000000000100000000011100010000000000000101000000000") port map( O =>C_0_S_3_L_6_out, I0 =>  inp_feat(282), I1 =>  inp_feat(85), I2 =>  inp_feat(249), I3 =>  inp_feat(255), I4 =>  inp_feat(15), I5 =>  inp_feat(323), I6 =>  inp_feat(94), I7 =>  inp_feat(345)); 
C_0_S_3_L_7_inst : LUT8 generic map(INIT => "0010101010100000000000000010000011100000101000000010100010100000101000101000000010100000000000001010000000000000000000000000000010001010100000000010101010101010110010001110000010101000111010100000000000000000000000100010100010100000000000000010000000100010") port map( O =>C_0_S_3_L_7_out, I0 =>  inp_feat(70), I1 =>  inp_feat(0), I2 =>  inp_feat(451), I3 =>  inp_feat(424), I4 =>  inp_feat(338), I5 =>  inp_feat(293), I6 =>  inp_feat(211), I7 =>  inp_feat(351)); 
C_0_S_4_L_0_inst : LUT8 generic map(INIT => "1111111011101110101011100000000001110000000000001010000000110000000011000100000010101010010000000000000000000000000000000000000011101110000001001010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_0_S_4_L_0_out, I0 =>  inp_feat(446), I1 =>  inp_feat(110), I2 =>  inp_feat(509), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_0_S_4_L_1_inst : LUT8 generic map(INIT => "0011000011100000101100001000000010111000110010001011000010100000101000101110101010000000001000001010000011000000000000000000000010101010100010001000000010000000100010001000100010000000100000001010000010000000100000000000000010100000100000000000000000000000") port map( O =>C_0_S_4_L_1_out, I0 =>  inp_feat(498), I1 =>  inp_feat(446), I2 =>  inp_feat(508), I3 =>  inp_feat(293), I4 =>  inp_feat(169), I5 =>  inp_feat(71), I6 =>  inp_feat(72), I7 =>  inp_feat(15)); 
C_0_S_4_L_2_inst : LUT8 generic map(INIT => "0011110111111101111111011100100011110111101100000111011111100000111000001100010011101100000000001000000010000000000000000000000011011100010100001000000000000000110000000000000001000000100000001000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_0_S_4_L_2_out, I0 =>  inp_feat(293), I1 =>  inp_feat(94), I2 =>  inp_feat(374), I3 =>  inp_feat(161), I4 =>  inp_feat(41), I5 =>  inp_feat(496), I6 =>  inp_feat(360), I7 =>  inp_feat(348)); 
C_0_S_4_L_3_inst : LUT8 generic map(INIT => "0101110011111100000000000000000011110000111110100000000000000000110011001110100010001000000000001000000011000000000000000000000011111101111111110000001000000000111000001011000000000000000000001110000000100000000000000000000011000000001000000000000000000000") port map( O =>C_0_S_4_L_3_out, I0 =>  inp_feat(41), I1 =>  inp_feat(319), I2 =>  inp_feat(259), I3 =>  inp_feat(222), I4 =>  inp_feat(70), I5 =>  inp_feat(61), I6 =>  inp_feat(111), I7 =>  inp_feat(249)); 
C_0_S_4_L_4_inst : LUT8 generic map(INIT => "1101110100001000000000000000000011111111000000001101000000000000110110100000000000000000000000001111100100000000000000000000000011111111110010001000000000000000111110010000000011110010000000001111010100000000000000000000000011111101000000000000000000000000") port map( O =>C_0_S_4_L_4_out, I0 =>  inp_feat(451), I1 =>  inp_feat(282), I2 =>  inp_feat(293), I3 =>  inp_feat(422), I4 =>  inp_feat(193), I5 =>  inp_feat(9), I6 =>  inp_feat(392), I7 =>  inp_feat(329)); 
C_0_S_4_L_5_inst : LUT8 generic map(INIT => "0110100010001000001011000000100000001000100010001000110010001000110010001000000010001000100000001000000010000000000000001000000010111011100000001111110110000000100010110000000000000000000000001000100010000000100010000000000000000000000000000000000000000000") port map( O =>C_0_S_4_L_5_out, I0 =>  inp_feat(42), I1 =>  inp_feat(485), I2 =>  inp_feat(9), I3 =>  inp_feat(496), I4 =>  inp_feat(338), I5 =>  inp_feat(347), I6 =>  inp_feat(293), I7 =>  inp_feat(329)); 
C_0_S_4_L_6_inst : LUT8 generic map(INIT => "1101100011111101100010001000000011011110111010001010100000001000011000001000000000000000000000001111110100101000101010000000100000000000111010000000100000000000101010001010100000000000000000001010000010100000000000000000000010100000101010000000100000001000") port map( O =>C_0_S_4_L_6_out, I0 =>  inp_feat(427), I1 =>  inp_feat(85), I2 =>  inp_feat(378), I3 =>  inp_feat(467), I4 =>  inp_feat(392), I5 =>  inp_feat(327), I6 =>  inp_feat(350), I7 =>  inp_feat(491)); 
C_0_S_4_L_7_inst : LUT8 generic map(INIT => "1110001011101111001100100010001111111110111011001111111000000000111001001110111000000000000000001100000011000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000011100100000000000000000010000000100010000000000000000000") port map( O =>C_0_S_4_L_7_out, I0 =>  inp_feat(338), I1 =>  inp_feat(72), I2 =>  inp_feat(130), I3 =>  inp_feat(302), I4 =>  inp_feat(379), I5 =>  inp_feat(71), I6 =>  inp_feat(9), I7 =>  inp_feat(193)); 
C_1_S_0_L_0_inst : LUT8 generic map(INIT => "1111101010001010100010000000000010101010101000101000101000000000100000001000000000000000000000000000000000000000000000000000000010101010000000101000110000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_1_S_0_L_0_out, I0 =>  inp_feat(463), I1 =>  inp_feat(287), I2 =>  inp_feat(480), I3 =>  inp_feat(42), I4 =>  inp_feat(358), I5 =>  inp_feat(462), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_1_S_0_L_1_inst : LUT8 generic map(INIT => "0001111110101000001011110000101001000010000000001100010000000000110011111000100000100010100010000000001100000000000000000000000011011111101010101100111110001110100011110000000011001111000000000000101000001010000011000000000000000000000000000000000000000000") port map( O =>C_1_S_0_L_1_out, I0 =>  inp_feat(74), I1 =>  inp_feat(439), I2 =>  inp_feat(293), I3 =>  inp_feat(72), I4 =>  inp_feat(88), I5 =>  inp_feat(59), I6 =>  inp_feat(110), I7 =>  inp_feat(328)); 
C_1_S_0_L_2_inst : LUT8 generic map(INIT => "0111011111111101111000001111100011000000110010000000000011000000111100001100000011100000110010000010000010101000100000001100100000000000000000000000000000001000000000001100000000000000000000001000100010001000100010001000100010001000100000001000100010001000") port map( O =>C_1_S_0_L_2_out, I0 =>  inp_feat(88), I1 =>  inp_feat(383), I2 =>  inp_feat(282), I3 =>  inp_feat(323), I4 =>  inp_feat(15), I5 =>  inp_feat(79), I6 =>  inp_feat(478), I7 =>  inp_feat(508)); 
C_1_S_0_L_3_inst : LUT8 generic map(INIT => "0111111111110100000000001101100011111010110100100000001001110000101010001010000010100000101010001011101110011011001000101011101000000000000000000000000000000000001111110000000000000010110010000000000010000000000000000000100000111011001110111010001010101010") port map( O =>C_1_S_0_L_3_out, I0 =>  inp_feat(293), I1 =>  inp_feat(478), I2 =>  inp_feat(289), I3 =>  inp_feat(272), I4 =>  inp_feat(390), I5 =>  inp_feat(180), I6 =>  inp_feat(302), I7 =>  inp_feat(282)); 
C_1_S_0_L_4_inst : LUT8 generic map(INIT => "1010111110101011101010001010100000001000000000001000100010001000101010101010101010101000101010001010100000000000101010001010000000000000000000000000000000000000000000000000000000001000000000001010000010100010000010000000000010101000000000001010100000000000") port map( O =>C_1_S_0_L_4_out, I0 =>  inp_feat(70), I1 =>  inp_feat(303), I2 =>  inp_feat(110), I3 =>  inp_feat(238), I4 =>  inp_feat(451), I5 =>  inp_feat(282), I6 =>  inp_feat(106), I7 =>  inp_feat(42)); 
C_1_S_0_L_5_inst : LUT8 generic map(INIT => "0010100100000111101000001110110011101010000000000100000010000000101111110000101100000000000000001010101000010000000000000100000010101010100010111010000011101110001010100000000011100000111000000011101101010011000000000010000110101010111000001110000011110000") port map( O =>C_1_S_0_L_5_out, I0 =>  inp_feat(483), I1 =>  inp_feat(302), I2 =>  inp_feat(180), I3 =>  inp_feat(6), I4 =>  inp_feat(496), I5 =>  inp_feat(121), I6 =>  inp_feat(329), I7 =>  inp_feat(212)); 
C_1_S_0_L_6_inst : LUT8 generic map(INIT => "0111001000100010101110100010001011101000000000001011100000101000110000010000000000100000000000001010100000000000101010001000100010110111001100000010000000000000101100000000000000000000001000001111111100100000101000000010000010100000000000001010000010100000") port map( O =>C_1_S_0_L_6_out, I0 =>  inp_feat(276), I1 =>  inp_feat(492), I2 =>  inp_feat(385), I3 =>  inp_feat(127), I4 =>  inp_feat(480), I5 =>  inp_feat(71), I6 =>  inp_feat(323), I7 =>  inp_feat(386)); 
C_1_S_0_L_7_inst : LUT8 generic map(INIT => "0100110000001100111011000000000010001100100000001110110110000000111111101010000010110000100000001000100010001000100000001000000011001100000000001000110000000000100010000000000001000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_1_S_0_L_7_out, I0 =>  inp_feat(480), I1 =>  inp_feat(337), I2 =>  inp_feat(452), I3 =>  inp_feat(292), I4 =>  inp_feat(323), I5 =>  inp_feat(381), I6 =>  inp_feat(446), I7 =>  inp_feat(360)); 
C_1_S_1_L_0_inst : LUT8 generic map(INIT => "1111101010001010100010000000000010101010101000101000101000000000100000001000000000000000000000000000000000000000000000000000000010101010000000101000110000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_1_S_1_L_0_out, I0 =>  inp_feat(463), I1 =>  inp_feat(287), I2 =>  inp_feat(480), I3 =>  inp_feat(42), I4 =>  inp_feat(358), I5 =>  inp_feat(462), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_1_S_1_L_1_inst : LUT8 generic map(INIT => "0010001110001110110011000000110010001110100000011100010011001100001110111000100010001000100010001111101110000000100000001000000010101010101011101010111000100100000000000000010001000100000001000000000000100000001000000010000000000000000000000000000000000000") port map( O =>C_1_S_1_L_1_out, I0 =>  inp_feat(462), I1 =>  inp_feat(351), I2 =>  inp_feat(468), I3 =>  inp_feat(166), I4 =>  inp_feat(72), I5 =>  inp_feat(129), I6 =>  inp_feat(110), I7 =>  inp_feat(328)); 
C_1_S_1_L_2_inst : LUT8 generic map(INIT => "0010111111111111101110101010001011100110101011111010001000000000000010101010101000001000001000101000100010100010000000000000000011101111111111111010101011111110111011110000111000000000000000001000101010001010001010100000101010001000000010000000000000000000") port map( O =>C_1_S_1_L_2_out, I0 =>  inp_feat(435), I1 =>  inp_feat(71), I2 =>  inp_feat(222), I3 =>  inp_feat(329), I4 =>  inp_feat(293), I5 =>  inp_feat(5), I6 =>  inp_feat(282), I7 =>  inp_feat(15)); 
C_1_S_1_L_3_inst : LUT8 generic map(INIT => "1111001011110000011000001111000010100000000000000000000000000000111100001110000011100000101000001111000010000000010000000000000000010000100000000000000000000000000100001000000000000000000000000001000010000000000000000000000010110000100000000000000000000000") port map( O =>C_1_S_1_L_3_out, I0 =>  inp_feat(169), I1 =>  inp_feat(90), I2 =>  inp_feat(70), I3 =>  inp_feat(61), I4 =>  inp_feat(402), I5 =>  inp_feat(261), I6 =>  inp_feat(302), I7 =>  inp_feat(282)); 
C_1_S_1_L_4_inst : LUT8 generic map(INIT => "1101100011011000100110001001100000001000000000001000100011001000000010001111100011111001111110001000000010000000000000001000100000011010100000001011101010001000000010001000000010001000100010001000101011001000101111111000100000000000100010001000001010001000") port map( O =>C_1_S_1_L_4_out, I0 =>  inp_feat(24), I1 =>  inp_feat(486), I2 =>  inp_feat(293), I3 =>  inp_feat(15), I4 =>  inp_feat(289), I5 =>  inp_feat(282), I6 =>  inp_feat(323), I7 =>  inp_feat(79)); 
C_1_S_1_L_5_inst : LUT8 generic map(INIT => "0000110000001000100010000000100011111100000001001000110000010100110010000000000010001000000010001000100000000000000011101000111111001110110001001100111101000100110011011000010011001101000001010000000000000000000000100000000000000000000000000000000000000000") port map( O =>C_1_S_1_L_5_out, I0 =>  inp_feat(323), I1 =>  inp_feat(42), I2 =>  inp_feat(302), I3 =>  inp_feat(390), I4 =>  inp_feat(9), I5 =>  inp_feat(108), I6 =>  inp_feat(446), I7 =>  inp_feat(249)); 
C_1_S_1_L_6_inst : LUT8 generic map(INIT => "0011001011110010101010101111001010110000101100101010000010101010111110101100101011000000110000000000000000000000000000000000000011101111110100111010100000000000101100010001000110100000000000001011001000000010000000000000000000100000000000000000000000000000") port map( O =>C_1_S_1_L_6_out, I0 =>  inp_feat(287), I1 =>  inp_feat(323), I2 =>  inp_feat(379), I3 =>  inp_feat(387), I4 =>  inp_feat(360), I5 =>  inp_feat(280), I6 =>  inp_feat(496), I7 =>  inp_feat(293)); 
C_1_S_1_L_7_inst : LUT8 generic map(INIT => "1000100001000000111011001101110011001000100000001100110011111111110101110101111110000000010000101100100000000000110001000100100011001000100000001100110011010100010010000011001001001000111111111110111011110010010000000001000010000000000000100100000011101000") port map( O =>C_1_S_1_L_7_out, I0 =>  inp_feat(372), I1 =>  inp_feat(508), I2 =>  inp_feat(484), I3 =>  inp_feat(287), I4 =>  inp_feat(427), I5 =>  inp_feat(450), I6 =>  inp_feat(265), I7 =>  inp_feat(272)); 
C_1_S_2_L_0_inst : LUT8 generic map(INIT => "1111101010001010100010000000000010101010101000101000101000000000100000001000000000000000000000000000000000000000000000000000000010101010000000101000110000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_1_S_2_L_0_out, I0 =>  inp_feat(463), I1 =>  inp_feat(287), I2 =>  inp_feat(480), I3 =>  inp_feat(42), I4 =>  inp_feat(358), I5 =>  inp_feat(462), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_1_S_2_L_1_inst : LUT8 generic map(INIT => "0010001110001110110011000000110010001110100000011100010011001100001110111000100010001000100010001111101110000000100000001000000010101010101011101010111000100100000000000000010001000100000001000000000000100000001000000010000000000000000000000000000000000000") port map( O =>C_1_S_2_L_1_out, I0 =>  inp_feat(462), I1 =>  inp_feat(351), I2 =>  inp_feat(468), I3 =>  inp_feat(166), I4 =>  inp_feat(72), I5 =>  inp_feat(129), I6 =>  inp_feat(110), I7 =>  inp_feat(328)); 
C_1_S_2_L_2_inst : LUT8 generic map(INIT => "0110111011101111101110101010001010101011101010100111000100000000000010100010101000001000001000101000100010100010000000000000000011101010111111111010101011101110101010100000100100000000000000001000101010001010001010100000101010001000000010000000000000000000") port map( O =>C_1_S_2_L_2_out, I0 =>  inp_feat(352), I1 =>  inp_feat(71), I2 =>  inp_feat(222), I3 =>  inp_feat(329), I4 =>  inp_feat(293), I5 =>  inp_feat(5), I6 =>  inp_feat(282), I7 =>  inp_feat(15)); 
C_1_S_2_L_3_inst : LUT8 generic map(INIT => "1101110011111101110000001111110111011100110101001100100011000100101100001111000000000000001100000001000001010100000000001100110001010000110000000000000000000000010100001101010000000000110010001101000000110000000000000000000001010000110100000000000011001100") port map( O =>C_1_S_2_L_3_out, I0 =>  inp_feat(308), I1 =>  inp_feat(319), I2 =>  inp_feat(275), I3 =>  inp_feat(108), I4 =>  inp_feat(53), I5 =>  inp_feat(9), I6 =>  inp_feat(451), I7 =>  inp_feat(282)); 
C_1_S_2_L_4_inst : LUT8 generic map(INIT => "1110110010110000111011001111010100000000010000001100000001000000101010001010000010101010101010001000100000000000010000000000000000101000000100000000000000010000000000000000000000000000000000001010000000000000000000000000000010000000000000000000000000000000") port map( O =>C_1_S_2_L_4_out, I0 =>  inp_feat(462), I1 =>  inp_feat(98), I2 =>  inp_feat(152), I3 =>  inp_feat(7), I4 =>  inp_feat(301), I5 =>  inp_feat(282), I6 =>  inp_feat(446), I7 =>  inp_feat(503)); 
C_1_S_2_L_5_inst : LUT8 generic map(INIT => "0001111001011101010011010101111111001000000010001100100000001000111010100000000011001000000000001100000000000000010000000000000011111110110110010000100010011001110010000000100011001000100010001010101000000000100000000000000011000000000000000000000000000000") port map( O =>C_1_S_2_L_5_out, I0 =>  inp_feat(58), I1 =>  inp_feat(485), I2 =>  inp_feat(222), I3 =>  inp_feat(451), I4 =>  inp_feat(331), I5 =>  inp_feat(293), I6 =>  inp_feat(360), I7 =>  inp_feat(323)); 
C_1_S_2_L_6_inst : LUT8 generic map(INIT => "1111100011100000011100001110000011100000101000001111000000010000111100001101000000110000101100001111000010100000011100000011000001110000011110000000000001000000000100001000000000000000000000001111000011010000000100001100000000010000000000000000000000000000") port map( O =>C_1_S_2_L_6_out, I0 =>  inp_feat(61), I1 =>  inp_feat(15), I2 =>  inp_feat(70), I3 =>  inp_feat(370), I4 =>  inp_feat(378), I5 =>  inp_feat(318), I6 =>  inp_feat(434), I7 =>  inp_feat(85)); 
C_1_S_2_L_7_inst : LUT8 generic map(INIT => "1000011001001000111011001100110001001110000000000010000000000000110011000000010011001100110001001000110000000000100000001000000010101010000010101011000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_1_S_2_L_7_out, I0 =>  inp_feat(348), I1 =>  inp_feat(219), I2 =>  inp_feat(293), I3 =>  inp_feat(390), I4 =>  inp_feat(302), I5 =>  inp_feat(275), I6 =>  inp_feat(153), I7 =>  inp_feat(288)); 
C_1_S_3_L_0_inst : LUT8 generic map(INIT => "1111101010001010100010000000000010101010101000101000101000000000100000001000000000000000000000000000000000000000000000000000000010101010000000101000110000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_1_S_3_L_0_out, I0 =>  inp_feat(463), I1 =>  inp_feat(287), I2 =>  inp_feat(480), I3 =>  inp_feat(42), I4 =>  inp_feat(358), I5 =>  inp_feat(462), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_1_S_3_L_1_inst : LUT8 generic map(INIT => "0000010011101100110011001100000011001100111011101000000000000000110011001000100011001100000000001100110010000000110011000000000000001100101000001010000000000000100010001110100011101010000000001000110010001000100001000000000010001000000000001000100000000000") port map( O =>C_1_S_3_L_1_out, I0 =>  inp_feat(323), I1 =>  inp_feat(498), I2 =>  inp_feat(509), I3 =>  inp_feat(446), I4 =>  inp_feat(288), I5 =>  inp_feat(71), I6 =>  inp_feat(15), I7 =>  inp_feat(328)); 
C_1_S_3_L_2_inst : LUT8 generic map(INIT => "0100110011001100000011000100000010001110110010000101010011110000110011001000000011001100000000000000010000000000010001000100000011000100110011001000000000000000100011000100010010000000000000001100100001000000110010000000000010000000000000000000000000000000") port map( O =>C_1_S_3_L_2_out, I0 =>  inp_feat(129), I1 =>  inp_feat(70), I2 =>  inp_feat(317), I3 =>  inp_feat(229), I4 =>  inp_feat(287), I5 =>  inp_feat(293), I6 =>  inp_feat(451), I7 =>  inp_feat(496)); 
C_1_S_3_L_3_inst : LUT8 generic map(INIT => "0010000010101110101000001000000010100000101010001010011010100000101011001100111110100000000000001010100010001000101000000000000000000100100010001100010000000000100000001000110011001100100000001000010010001100100001000000000010001100100011001000010000000000") port map( O =>C_1_S_3_L_3_out, I0 =>  inp_feat(499), I1 =>  inp_feat(360), I2 =>  inp_feat(386), I3 =>  inp_feat(478), I4 =>  inp_feat(241), I5 =>  inp_feat(41), I6 =>  inp_feat(222), I7 =>  inp_feat(468)); 
C_1_S_3_L_4_inst : LUT8 generic map(INIT => "1111110111100000100010001010000010101000101011000000000000101100000000000000000010100000000000001010100010101100001000100010100001000000110001001101000011010000000010000000110000000000000011000010000000100000000000000000000000000000101010000000000000101010") port map( O =>C_1_S_3_L_4_out, I0 =>  inp_feat(99), I1 =>  inp_feat(388), I2 =>  inp_feat(172), I3 =>  inp_feat(376), I4 =>  inp_feat(390), I5 =>  inp_feat(381), I6 =>  inp_feat(287), I7 =>  inp_feat(436)); 
C_1_S_3_L_5_inst : LUT8 generic map(INIT => "0101101111001010101010101000110000001010101010100000000000000000111101001101000011110000110110000000000010000000000000001000000011011111110011000000100011001100000000000000000000000000000000001100110001001000000000001100100000000000000000000000000000000000") port map( O =>C_1_S_3_L_5_out, I0 =>  inp_feat(317), I1 =>  inp_feat(390), I2 =>  inp_feat(222), I3 =>  inp_feat(72), I4 =>  inp_feat(166), I5 =>  inp_feat(258), I6 =>  inp_feat(293), I7 =>  inp_feat(506)); 
C_1_S_3_L_6_inst : LUT8 generic map(INIT => "1100100010110000111100001111010010000000001000001011010011110000000000000011000000000000110100000000000000000000000100000000000010001000000000001001100000010000100010000000000000000000000000000000100000110000000110000011000000000000000000000100000000000000") port map( O =>C_1_S_3_L_6_out, I0 =>  inp_feat(348), I1 =>  inp_feat(338), I2 =>  inp_feat(59), I3 =>  inp_feat(110), I4 =>  inp_feat(323), I5 =>  inp_feat(47), I6 =>  inp_feat(282), I7 =>  inp_feat(9)); 
C_1_S_3_L_7_inst : LUT8 generic map(INIT => "1110111110001100110111111100010011101010110010001100001000000000110000001100000001000000000000001110100011100000000000000000000001101000010000001100000000000000100010100000100000000000000000001100100001000000100000000000000010000000000000000000000000000000") port map( O =>C_1_S_3_L_7_out, I0 =>  inp_feat(293), I1 =>  inp_feat(359), I2 =>  inp_feat(388), I3 =>  inp_feat(440), I4 =>  inp_feat(436), I5 =>  inp_feat(339), I6 =>  inp_feat(411), I7 =>  inp_feat(170)); 
C_1_S_4_L_0_inst : LUT8 generic map(INIT => "1111101010001010100010000000000010101010101000101000101000000000100000001000000000000000000000000000000000000000000000000000000010101010000000101000110000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_1_S_4_L_0_out, I0 =>  inp_feat(463), I1 =>  inp_feat(287), I2 =>  inp_feat(480), I3 =>  inp_feat(42), I4 =>  inp_feat(358), I5 =>  inp_feat(462), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_1_S_4_L_1_inst : LUT8 generic map(INIT => "0100110000000000110010000000000011001110000010001000100010000000110011001000100011000000000000001100110000000000110000000000000010001100000000001010000010000000110011001000100010001000100010001100110010001000100001001000000010001100000000001000010010000000") port map( O =>C_1_S_4_L_1_out, I0 =>  inp_feat(212), I1 =>  inp_feat(70), I2 =>  inp_feat(310), I3 =>  inp_feat(173), I4 =>  inp_feat(288), I5 =>  inp_feat(71), I6 =>  inp_feat(15), I7 =>  inp_feat(328)); 
C_1_S_4_L_2_inst : LUT8 generic map(INIT => "1000011000000000101011100000000000000000000010000000100010001000111111110000000011101010000000000000100000000000100010000000100011101110110001001100111001001110110000001100000010100000000000001100000000000000100000000000000010000000000000001000000000000000") port map( O =>C_1_S_4_L_2_out, I0 =>  inp_feat(350), I1 =>  inp_feat(318), I2 =>  inp_feat(75), I3 =>  inp_feat(42), I4 =>  inp_feat(108), I5 =>  inp_feat(287), I6 =>  inp_feat(293), I7 =>  inp_feat(302)); 
C_1_S_4_L_3_inst : LUT8 generic map(INIT => "1110110001111111110011000101111100000000000000001110000010000000111100101011111111110000101010100111000010100000111100001010000001100000001001110100000000000000000000000000000000000000000000001111000000101111000000000000000001000000000000100000000000000000") port map( O =>C_1_S_4_L_3_out, I0 =>  inp_feat(71), I1 =>  inp_feat(222), I2 =>  inp_feat(10), I3 =>  inp_feat(245), I4 =>  inp_feat(75), I5 =>  inp_feat(485), I6 =>  inp_feat(302), I7 =>  inp_feat(287)); 
C_1_S_4_L_4_inst : LUT8 generic map(INIT => "0111111111111000000100001010101010110001101100000010000110100000110000000000000000001110000000100000000000000000101011101010001000111111110011000000000000000000001100000010000000000000000000000000010000000000000001110000000000000000000000001010111000000000") port map( O =>C_1_S_4_L_4_out, I0 =>  inp_feat(61), I1 =>  inp_feat(297), I2 =>  inp_feat(380), I3 =>  inp_feat(350), I4 =>  inp_feat(338), I5 =>  inp_feat(110), I6 =>  inp_feat(237), I7 =>  inp_feat(378)); 
C_1_S_4_L_5_inst : LUT8 generic map(INIT => "1101111011110000100000101000101000000000100000001010001010000010000000000101000000000000001000000000000000000000001000000010001011111010001100001000000000000000001100100011001000100010001100100011000000000000000000100000000000000000000000100010001000100010") port map( O =>C_1_S_4_L_5_out, I0 =>  inp_feat(470), I1 =>  inp_feat(172), I2 =>  inp_feat(462), I3 =>  inp_feat(110), I4 =>  inp_feat(348), I5 =>  inp_feat(338), I6 =>  inp_feat(282), I7 =>  inp_feat(302)); 
C_1_S_4_L_6_inst : LUT8 generic map(INIT => "1010111000001110101110110011110100001100001010000010001100110001100010000000100010110001001100001000100010000000101100011011001100101100000010001010000010001100000000000000000000000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_1_S_4_L_6_out, I0 =>  inp_feat(508), I1 =>  inp_feat(338), I2 =>  inp_feat(293), I3 =>  inp_feat(33), I4 =>  inp_feat(308), I5 =>  inp_feat(282), I6 =>  inp_feat(9), I7 =>  inp_feat(275)); 
C_1_S_4_L_7_inst : LUT8 generic map(INIT => "0010011110000010000000101111101101000010100000100110101011111011111011101000000000000000100010000000100010000000100010001000100011111010110000000000000011000000100000001100000000000000110000001110111011000000000000000100000001000000110000000000000001000000") port map( O =>C_1_S_4_L_7_out, I0 =>  inp_feat(476), I1 =>  inp_feat(229), I2 =>  inp_feat(303), I3 =>  inp_feat(293), I4 =>  inp_feat(224), I5 =>  inp_feat(493), I6 =>  inp_feat(327), I7 =>  inp_feat(415)); 
C_2_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000001000100010001000000000000000000000000000000010000000000000000000000010000000100000000000000000000000000010000000000000000000000010001000100010000000000000000000") port map( O =>C_2_S_0_L_0_out, I0 =>  inp_feat(327), I1 =>  inp_feat(297), I2 =>  inp_feat(155), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_2_S_0_L_1_inst : LUT8 generic map(INIT => "1110000110100010000000000000000000000000100000000000000000000000000000000011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_0_L_1_out, I0 =>  inp_feat(233), I1 =>  inp_feat(378), I2 =>  inp_feat(314), I3 =>  inp_feat(287), I4 =>  inp_feat(293), I5 =>  inp_feat(329), I6 =>  inp_feat(241), I7 =>  inp_feat(478)); 
C_2_S_0_L_2_inst : LUT8 generic map(INIT => "1100000000000000000000000000000011010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_0_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(386), I2 =>  inp_feat(446), I3 =>  inp_feat(211), I4 =>  inp_feat(71), I5 =>  inp_feat(465), I6 =>  inp_feat(351), I7 =>  inp_feat(72)); 
C_2_S_0_L_3_inst : LUT8 generic map(INIT => "0100100000000000000001000000000000000000000000001100010000000000000000000000000000000000000000001000000000000000100000000000000010001100000001000000000000000000000010010000000001000100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_0_L_3_out, I0 =>  inp_feat(42), I1 =>  inp_feat(106), I2 =>  inp_feat(282), I3 =>  inp_feat(90), I4 =>  inp_feat(70), I5 =>  inp_feat(462), I6 =>  inp_feat(477), I7 =>  inp_feat(193)); 
C_2_S_0_L_4_inst : LUT8 generic map(INIT => "0000100000000000100010000000000000000000000000000000000000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_0_L_4_out, I0 =>  inp_feat(374), I1 =>  inp_feat(450), I2 =>  inp_feat(439), I3 =>  inp_feat(24), I4 =>  inp_feat(122), I5 =>  inp_feat(348), I6 =>  inp_feat(440), I7 =>  inp_feat(327)); 
C_2_S_0_L_5_inst : LUT8 generic map(INIT => "0110100000000000000000000000000000101010000000000000000000000000000000000000000000000000000000001010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000") port map( O =>C_2_S_0_L_5_out, I0 =>  inp_feat(40), I1 =>  inp_feat(127), I2 =>  inp_feat(355), I3 =>  inp_feat(505), I4 =>  inp_feat(478), I5 =>  inp_feat(462), I6 =>  inp_feat(215), I7 =>  inp_feat(71)); 
C_2_S_0_L_6_inst : LUT8 generic map(INIT => "0010000000000000000000000000000010101000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000101000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000") port map( O =>C_2_S_0_L_6_out, I0 =>  inp_feat(348), I1 =>  inp_feat(347), I2 =>  inp_feat(509), I3 =>  inp_feat(293), I4 =>  inp_feat(306), I5 =>  inp_feat(127), I6 =>  inp_feat(95), I7 =>  inp_feat(85)); 
C_2_S_0_L_7_inst : LUT8 generic map(INIT => "0010110010101010000010001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_0_L_7_out, I0 =>  inp_feat(318), I1 =>  inp_feat(355), I2 =>  inp_feat(345), I3 =>  inp_feat(215), I4 =>  inp_feat(323), I5 =>  inp_feat(370), I6 =>  inp_feat(219), I7 =>  inp_feat(90)); 
C_2_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000001000100010001000000000000000000000000000000010000000000000000000000010000000100000000000000000000000000010000000000000000000000010001000100010000000000000000000") port map( O =>C_2_S_1_L_0_out, I0 =>  inp_feat(327), I1 =>  inp_feat(297), I2 =>  inp_feat(155), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_2_S_1_L_1_inst : LUT8 generic map(INIT => "1110000110100010000000000000000000000000100000000000000000000000000000000011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_1_L_1_out, I0 =>  inp_feat(233), I1 =>  inp_feat(378), I2 =>  inp_feat(314), I3 =>  inp_feat(287), I4 =>  inp_feat(293), I5 =>  inp_feat(329), I6 =>  inp_feat(241), I7 =>  inp_feat(478)); 
C_2_S_1_L_2_inst : LUT8 generic map(INIT => "1100000000000000000000000000000011010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_1_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(386), I2 =>  inp_feat(446), I3 =>  inp_feat(211), I4 =>  inp_feat(71), I5 =>  inp_feat(465), I6 =>  inp_feat(351), I7 =>  inp_feat(72)); 
C_2_S_1_L_3_inst : LUT8 generic map(INIT => "0000001000001000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010000000001010101000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_1_L_3_out, I0 =>  inp_feat(75), I1 =>  inp_feat(260), I2 =>  inp_feat(130), I3 =>  inp_feat(62), I4 =>  inp_feat(192), I5 =>  inp_feat(348), I6 =>  inp_feat(327), I7 =>  inp_feat(282)); 
C_2_S_1_L_4_inst : LUT8 generic map(INIT => "0110110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_1_L_4_out, I0 =>  inp_feat(177), I1 =>  inp_feat(376), I2 =>  inp_feat(287), I3 =>  inp_feat(71), I4 =>  inp_feat(478), I5 =>  inp_feat(348), I6 =>  inp_feat(327), I7 =>  inp_feat(282)); 
C_2_S_1_L_5_inst : LUT8 generic map(INIT => "0001000000000000111100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000001111000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_1_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(396), I2 =>  inp_feat(68), I3 =>  inp_feat(108), I4 =>  inp_feat(440), I5 =>  inp_feat(88), I6 =>  inp_feat(371), I7 =>  inp_feat(193)); 
C_2_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000001000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_1_L_6_out, I0 =>  inp_feat(269), I1 =>  inp_feat(327), I2 =>  inp_feat(348), I3 =>  inp_feat(446), I4 =>  inp_feat(178), I5 =>  inp_feat(440), I6 =>  inp_feat(415), I7 =>  inp_feat(122)); 
C_2_S_1_L_7_inst : LUT8 generic map(INIT => "1010100000000000101000001000000000000000001000001010000010100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000") port map( O =>C_2_S_1_L_7_out, I0 =>  inp_feat(293), I1 =>  inp_feat(440), I2 =>  inp_feat(302), I3 =>  inp_feat(193), I4 =>  inp_feat(465), I5 =>  inp_feat(82), I6 =>  inp_feat(478), I7 =>  inp_feat(323)); 
C_2_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000001000100010001000000000000000000000000000000010000000000000000000000010000000100000000000000000000000000010000000000000000000000010001000100010000000000000000000") port map( O =>C_2_S_2_L_0_out, I0 =>  inp_feat(327), I1 =>  inp_feat(297), I2 =>  inp_feat(155), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_2_S_2_L_1_inst : LUT8 generic map(INIT => "1111000001010000110000000000000000000000000000000001000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_2_L_1_out, I0 =>  inp_feat(282), I1 =>  inp_feat(504), I2 =>  inp_feat(327), I3 =>  inp_feat(442), I4 =>  inp_feat(287), I5 =>  inp_feat(329), I6 =>  inp_feat(241), I7 =>  inp_feat(478)); 
C_2_S_2_L_2_inst : LUT8 generic map(INIT => "1010001000000010101000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_2_L_2_out, I0 =>  inp_feat(293), I1 =>  inp_feat(155), I2 =>  inp_feat(329), I3 =>  inp_feat(226), I4 =>  inp_feat(465), I5 =>  inp_feat(245), I6 =>  inp_feat(71), I7 =>  inp_feat(72)); 
C_2_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000100000000000000000000000100000001000000000000000000000000000000010000000000000000000000000000000100010000000000000000000000000001000100000000000000000000000000010001000000000000000000000000000") port map( O =>C_2_S_2_L_3_out, I0 =>  inp_feat(446), I1 =>  inp_feat(348), I2 =>  inp_feat(139), I3 =>  inp_feat(41), I4 =>  inp_feat(99), I5 =>  inp_feat(401), I6 =>  inp_feat(152), I7 =>  inp_feat(440)); 
C_2_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000010101000000000000010100000000000001010000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_2_L_4_out, I0 =>  inp_feat(222), I1 =>  inp_feat(379), I2 =>  inp_feat(289), I3 =>  inp_feat(108), I4 =>  inp_feat(347), I5 =>  inp_feat(462), I6 =>  inp_feat(37), I7 =>  inp_feat(478)); 
C_2_S_2_L_5_inst : LUT8 generic map(INIT => "0000100000001000100010000000100010101000000000001000100000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_2_L_5_out, I0 =>  inp_feat(386), I1 =>  inp_feat(75), I2 =>  inp_feat(42), I3 =>  inp_feat(108), I4 =>  inp_feat(347), I5 =>  inp_feat(462), I6 =>  inp_feat(37), I7 =>  inp_feat(478)); 
C_2_S_2_L_6_inst : LUT8 generic map(INIT => "0010000000000000000000000000000010100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000101000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_2_L_6_out, I0 =>  inp_feat(5), I1 =>  inp_feat(388), I2 =>  inp_feat(71), I3 =>  inp_feat(222), I4 =>  inp_feat(323), I5 =>  inp_feat(378), I6 =>  inp_feat(452), I7 =>  inp_feat(215)); 
C_2_S_2_L_7_inst : LUT8 generic map(INIT => "0010001000100000100000100000000000000000000000000000101000000000001000100000000000100010000000001000000000000000000000000000000000100000000000000010000000000000000000000000000000000000010000001010001000000000001000100100000000000000000000000000000000000000") port map( O =>C_2_S_2_L_7_out, I0 =>  inp_feat(68), I1 =>  inp_feat(70), I2 =>  inp_feat(83), I3 =>  inp_feat(323), I4 =>  inp_feat(190), I5 =>  inp_feat(391), I6 =>  inp_feat(193), I7 =>  inp_feat(206)); 
C_2_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000001000100010001000000000000000000000000000000010000000000000000000000010000000100000000000000000000000000010000000000000000000000010001000100010000000000000000000") port map( O =>C_2_S_3_L_0_out, I0 =>  inp_feat(327), I1 =>  inp_feat(297), I2 =>  inp_feat(155), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_2_S_3_L_1_inst : LUT8 generic map(INIT => "1111000001010000110000000000000000000000000000000001000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_1_out, I0 =>  inp_feat(282), I1 =>  inp_feat(504), I2 =>  inp_feat(327), I3 =>  inp_feat(442), I4 =>  inp_feat(287), I5 =>  inp_feat(329), I6 =>  inp_feat(241), I7 =>  inp_feat(478)); 
C_2_S_3_L_2_inst : LUT8 generic map(INIT => "1110000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_2_out, I0 =>  inp_feat(386), I1 =>  inp_feat(323), I2 =>  inp_feat(156), I3 =>  inp_feat(394), I4 =>  inp_feat(495), I5 =>  inp_feat(25), I6 =>  inp_feat(71), I7 =>  inp_feat(72)); 
C_2_S_3_L_3_inst : LUT8 generic map(INIT => "0000000010000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_3_out, I0 =>  inp_feat(496), I1 =>  inp_feat(75), I2 =>  inp_feat(41), I3 =>  inp_feat(401), I4 =>  inp_feat(152), I5 =>  inp_feat(348), I6 =>  inp_feat(92), I7 =>  inp_feat(440)); 
C_2_S_3_L_4_inst : LUT8 generic map(INIT => "0100110000000000000000000000000000001000000000000100000000000000110011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_4_out, I0 =>  inp_feat(358), I1 =>  inp_feat(293), I2 =>  inp_feat(345), I3 =>  inp_feat(72), I4 =>  inp_feat(386), I5 =>  inp_feat(509), I6 =>  inp_feat(347), I7 =>  inp_feat(327)); 
C_2_S_3_L_5_inst : LUT8 generic map(INIT => "0100000011101101000000000001000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000011011000111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_5_out, I0 =>  inp_feat(345), I1 =>  inp_feat(437), I2 =>  inp_feat(432), I3 =>  inp_feat(282), I4 =>  inp_feat(289), I5 =>  inp_feat(302), I6 =>  inp_feat(293), I7 =>  inp_feat(192)); 
C_2_S_3_L_6_inst : LUT8 generic map(INIT => "0000100000001000100000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_6_out, I0 =>  inp_feat(298), I1 =>  inp_feat(243), I2 =>  inp_feat(42), I3 =>  inp_feat(90), I4 =>  inp_feat(487), I5 =>  inp_feat(354), I6 =>  inp_feat(450), I7 =>  inp_feat(3)); 
C_2_S_3_L_7_inst : LUT8 generic map(INIT => "1100000010000000011100001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_3_L_7_out, I0 =>  inp_feat(195), I1 =>  inp_feat(48), I2 =>  inp_feat(348), I3 =>  inp_feat(42), I4 =>  inp_feat(357), I5 =>  inp_feat(289), I6 =>  inp_feat(293), I7 =>  inp_feat(302)); 
C_2_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000001000100010001000000000000000000000000000000010000000000000000000000010000000100000000000000000000000000010000000000000000000000010001000100010000000000000000000") port map( O =>C_2_S_4_L_0_out, I0 =>  inp_feat(327), I1 =>  inp_feat(297), I2 =>  inp_feat(155), I3 =>  inp_feat(485), I4 =>  inp_feat(33), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_2_S_4_L_1_inst : LUT8 generic map(INIT => "1111000001010000110000000000000000000000000000000001000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_4_L_1_out, I0 =>  inp_feat(282), I1 =>  inp_feat(504), I2 =>  inp_feat(327), I3 =>  inp_feat(442), I4 =>  inp_feat(287), I5 =>  inp_feat(329), I6 =>  inp_feat(241), I7 =>  inp_feat(478)); 
C_2_S_4_L_2_inst : LUT8 generic map(INIT => "1010000000000000100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_4_L_2_out, I0 =>  inp_feat(386), I1 =>  inp_feat(260), I2 =>  inp_feat(9), I3 =>  inp_feat(72), I4 =>  inp_feat(142), I5 =>  inp_feat(438), I6 =>  inp_feat(71), I7 =>  inp_feat(211)); 
C_2_S_4_L_3_inst : LUT8 generic map(INIT => "0010000000000000100000000000000000000000000000000000000000000000111000001000000011100000100000000000000000000000000000000000000010100000000100000000000100000000000000000000000000000000000100001010000000100000101000000000000000000000000000000000000000000000") port map( O =>C_2_S_4_L_3_out, I0 =>  inp_feat(323), I1 =>  inp_feat(357), I2 =>  inp_feat(222), I3 =>  inp_feat(134), I4 =>  inp_feat(390), I5 =>  inp_feat(71), I6 =>  inp_feat(192), I7 =>  inp_feat(190)); 
C_2_S_4_L_4_inst : LUT8 generic map(INIT => "1000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_4_L_4_out, I0 =>  inp_feat(293), I1 =>  inp_feat(90), I2 =>  inp_feat(348), I3 =>  inp_feat(219), I4 =>  inp_feat(72), I5 =>  inp_feat(41), I6 =>  inp_feat(509), I7 =>  inp_feat(178)); 
C_2_S_4_L_5_inst : LUT8 generic map(INIT => "0100000000000000110000000000000000000000000000000000000000000000110011000000000011001100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_4_L_5_out, I0 =>  inp_feat(485), I1 =>  inp_feat(348), I2 =>  inp_feat(197), I3 =>  inp_feat(211), I4 =>  inp_feat(432), I5 =>  inp_feat(441), I6 =>  inp_feat(440), I7 =>  inp_feat(327)); 
C_2_S_4_L_6_inst : LUT8 generic map(INIT => "0010000000000000100000000000000010000001000000001000000000000000000000000000000000000000000000001000000000000000000000000000000010100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_2_S_4_L_6_out, I0 =>  inp_feat(71), I1 =>  inp_feat(220), I2 =>  inp_feat(478), I3 =>  inp_feat(290), I4 =>  inp_feat(482), I5 =>  inp_feat(287), I6 =>  inp_feat(493), I7 =>  inp_feat(3)); 
C_2_S_4_L_7_inst : LUT8 generic map(INIT => "0100000000000000001000000000000001010101010101000111010101010000000000000001000000000000000000000001000000010000000000000000000000010000000001001000000000000000111100000101010011110000010100000000000000000000000000000000000000000000010000000000000000000000") port map( O =>C_2_S_4_L_7_out, I0 =>  inp_feat(413), I1 =>  inp_feat(378), I2 =>  inp_feat(62), I3 =>  inp_feat(149), I4 =>  inp_feat(486), I5 =>  inp_feat(508), I6 =>  inp_feat(323), I7 =>  inp_feat(379)); 
C_3_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000101000010000000000110000100100001010000000000000000000000000000011000000000000000010000000000000110010000000000000000000000000001000000000000000000000000000000010100000000000000000000000000000") port map( O =>C_3_S_0_L_0_out, I0 =>  inp_feat(220), I1 =>  inp_feat(210), I2 =>  inp_feat(372), I3 =>  inp_feat(340), I4 =>  inp_feat(90), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_3_S_0_L_1_inst : LUT8 generic map(INIT => "1011011011111010000000000000000000000000100000000000000000000000000000000110100000000000000000000000000000000000000000000000000011111110011100111000000100100111000000000000000000000000000000001111111111010000110000000000000000000000000000000000000000000000") port map( O =>C_3_S_0_L_1_out, I0 =>  inp_feat(83), I1 =>  inp_feat(331), I2 =>  inp_feat(201), I3 =>  inp_feat(504), I4 =>  inp_feat(327), I5 =>  inp_feat(50), I6 =>  inp_feat(340), I7 =>  inp_feat(337)); 
C_3_S_0_L_2_inst : LUT8 generic map(INIT => "1010000000000001000000000000000000100000000100010000000000000000000010000010000000000000000000001000100000000000000010000000000010001000000000000000000000000000101000000001000100000000000000000000100000000000000000000000000000101000000000000000100000000000") port map( O =>C_3_S_0_L_2_out, I0 =>  inp_feat(376), I1 =>  inp_feat(70), I2 =>  inp_feat(11), I3 =>  inp_feat(224), I4 =>  inp_feat(311), I5 =>  inp_feat(508), I6 =>  inp_feat(503), I7 =>  inp_feat(440)); 
C_3_S_0_L_3_inst : LUT8 generic map(INIT => "0101110001001000000000001110000001010000000000001101000000000000000000000000000000000000000000000000000000000000000000001000000010000000110000000000000011000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_0_L_3_out, I0 =>  inp_feat(355), I1 =>  inp_feat(71), I2 =>  inp_feat(461), I3 =>  inp_feat(152), I4 =>  inp_feat(77), I5 =>  inp_feat(224), I6 =>  inp_feat(143), I7 =>  inp_feat(503)); 
C_3_S_0_L_4_inst : LUT8 generic map(INIT => "1000001010011010000001000000000001110111010100010000000000000000111001011100110011001101110000001101111100101101010001000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_3_S_0_L_4_out, I0 =>  inp_feat(282), I1 =>  inp_feat(201), I2 =>  inp_feat(290), I3 =>  inp_feat(500), I4 =>  inp_feat(339), I5 =>  inp_feat(470), I6 =>  inp_feat(152), I7 =>  inp_feat(143)); 
C_3_S_0_L_5_inst : LUT8 generic map(INIT => "0110000000000000000100000000000010010000000000000000000000000000111101000100010101010001000100001000000000000000000000000000000011000000010001000000000001000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_0_L_5_out, I0 =>  inp_feat(285), I1 =>  inp_feat(499), I2 =>  inp_feat(445), I3 =>  inp_feat(296), I4 =>  inp_feat(242), I5 =>  inp_feat(467), I6 =>  inp_feat(465), I7 =>  inp_feat(77)); 
C_3_S_0_L_6_inst : LUT8 generic map(INIT => "1000101000101011101000000011101100000000000000000000000010000000100000001001011110000000010000111000000010000000100000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_0_L_6_out, I0 =>  inp_feat(277), I1 =>  inp_feat(70), I2 =>  inp_feat(192), I3 =>  inp_feat(65), I4 =>  inp_feat(149), I5 =>  inp_feat(116), I6 =>  inp_feat(83), I7 =>  inp_feat(143)); 
C_3_S_0_L_7_inst : LUT8 generic map(INIT => "1111101110100010000010100000001101100001000000000000000000000000000100000000000000000000000000011010000000000000000000000000000001011100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_0_L_7_out, I0 =>  inp_feat(154), I1 =>  inp_feat(282), I2 =>  inp_feat(295), I3 =>  inp_feat(432), I4 =>  inp_feat(461), I5 =>  inp_feat(201), I6 =>  inp_feat(327), I7 =>  inp_feat(41)); 
C_3_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000001000010000000000000000000000000000000000000000000000100011001010100000001001000000000000000000001011100000000000101111001000100010000000000000000000100000001100000001000100010001000000000000001100000000000000000000000000000000000000000000000000") port map( O =>C_3_S_1_L_0_out, I0 =>  inp_feat(259), I1 =>  inp_feat(340), I2 =>  inp_feat(82), I3 =>  inp_feat(83), I4 =>  inp_feat(161), I5 =>  inp_feat(141), I6 =>  inp_feat(483), I7 =>  inp_feat(421)); 
C_3_S_1_L_1_inst : LUT8 generic map(INIT => "1110000000110000100010000010000010100000011100000011000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_1_L_1_out, I0 =>  inp_feat(297), I1 =>  inp_feat(183), I2 =>  inp_feat(403), I3 =>  inp_feat(87), I4 =>  inp_feat(298), I5 =>  inp_feat(494), I6 =>  inp_feat(266), I7 =>  inp_feat(143)); 
C_3_S_1_L_2_inst : LUT8 generic map(INIT => "1000000011100000000000000000000000010000001000000000000000000000000000000000110000000000000000000000000000000000000000000000000000100011101000000000000000000000001000001010000000000000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_1_L_2_out, I0 =>  inp_feat(5), I1 =>  inp_feat(98), I2 =>  inp_feat(9), I3 =>  inp_feat(508), I4 =>  inp_feat(311), I5 =>  inp_feat(11), I6 =>  inp_feat(403), I7 =>  inp_feat(258)); 
C_3_S_1_L_3_inst : LUT8 generic map(INIT => "0100110000110000100000000000000000000000000000000000000000000000100001000000000010001100000001000000000000000000000011000000000000100010111100101000000000000000100010000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_3_S_1_L_3_out, I0 =>  inp_feat(492), I1 =>  inp_feat(391), I2 =>  inp_feat(427), I3 =>  inp_feat(442), I4 =>  inp_feat(465), I5 =>  inp_feat(296), I6 =>  inp_feat(402), I7 =>  inp_feat(440)); 
C_3_S_1_L_4_inst : LUT8 generic map(INIT => "1111100000100000101110000001000000100000000000100000001100000010111100000000000010100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000011000000001000000000001000100010001000000000000000000000000000001000000010") port map( O =>C_3_S_1_L_4_out, I0 =>  inp_feat(376), I1 =>  inp_feat(473), I2 =>  inp_feat(323), I3 =>  inp_feat(212), I4 =>  inp_feat(6), I5 =>  inp_feat(116), I6 =>  inp_feat(193), I7 =>  inp_feat(467)); 
C_3_S_1_L_5_inst : LUT8 generic map(INIT => "1100001100000101000000000000000000000000000010000010000000000000000000000001010000100000000000000000000000000000101010000000000011111100000000001100000000000000010000000000000000000000000000000100010000000000000000000000000100000000000000000000000000000000") port map( O =>C_3_S_1_L_5_out, I0 =>  inp_feat(209), I1 =>  inp_feat(483), I2 =>  inp_feat(468), I3 =>  inp_feat(374), I4 =>  inp_feat(503), I5 =>  inp_feat(148), I6 =>  inp_feat(93), I7 =>  inp_feat(70)); 
C_3_S_1_L_6_inst : LUT8 generic map(INIT => "0000010000000000000000000000000001000000000000000100000001000000000000000000000000010100010101001000000000000000010000000101010100100000100000000001010000000000000000000000000011011111000000000000000000000000000111100000000000000101000010000000110100001111") port map( O =>C_3_S_1_L_6_out, I0 =>  inp_feat(462), I1 =>  inp_feat(93), I2 =>  inp_feat(427), I3 =>  inp_feat(394), I4 =>  inp_feat(70), I5 =>  inp_feat(192), I6 =>  inp_feat(77), I7 =>  inp_feat(158)); 
C_3_S_1_L_7_inst : LUT8 generic map(INIT => "1101111001010000000000010000000001001100000000000100010100000101001111010100000010000001000000001100010100000000000000000000000000000001000001000000000100000000000001010000010000000101000000000000000000000000000000000100000100000000000000000000010001000000") port map( O =>C_3_S_1_L_7_out, I0 =>  inp_feat(282), I1 =>  inp_feat(467), I2 =>  inp_feat(152), I3 =>  inp_feat(327), I4 =>  inp_feat(259), I5 =>  inp_feat(83), I6 =>  inp_feat(65), I7 =>  inp_feat(328)); 
C_3_S_2_L_0_inst : LUT8 generic map(INIT => "1101100010001000000000000000000010101010001000000010000000000000000000000010000100000000000000000010001000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_2_L_0_out, I0 =>  inp_feat(11), I1 =>  inp_feat(232), I2 =>  inp_feat(281), I3 =>  inp_feat(77), I4 =>  inp_feat(266), I5 =>  inp_feat(209), I6 =>  inp_feat(494), I7 =>  inp_feat(143)); 
C_3_S_2_L_1_inst : LUT8 generic map(INIT => "0001000101000000110000000000000000000000000000011000100000000000111100010101100110100000000000000000000101011011000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000") port map( O =>C_3_S_2_L_1_out, I0 =>  inp_feat(508), I1 =>  inp_feat(442), I2 =>  inp_feat(386), I3 =>  inp_feat(400), I4 =>  inp_feat(468), I5 =>  inp_feat(493), I6 =>  inp_feat(347), I7 =>  inp_feat(311)); 
C_3_S_2_L_2_inst : LUT8 generic map(INIT => "1010000000000000001000000000000010000010000000010000000100000000001110100000000010000000000000001011101100000001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000100000000") port map( O =>C_3_S_2_L_2_out, I0 =>  inp_feat(166), I1 =>  inp_feat(198), I2 =>  inp_feat(400), I3 =>  inp_feat(458), I4 =>  inp_feat(37), I5 =>  inp_feat(258), I6 =>  inp_feat(508), I7 =>  inp_feat(311)); 
C_3_S_2_L_3_inst : LUT8 generic map(INIT => "1100001001001000000000001010100000000000000000000000000010100000110000001100000010000000100010000010000000100000100000001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000100000000000000000000000000010000000") port map( O =>C_3_S_2_L_3_out, I0 =>  inp_feat(427), I1 =>  inp_feat(212), I2 =>  inp_feat(458), I3 =>  inp_feat(347), I4 =>  inp_feat(258), I5 =>  inp_feat(110), I6 =>  inp_feat(508), I7 =>  inp_feat(311)); 
C_3_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000001000010001000000000100010000100011000000000000000000000000000000100100000000000000001000000000000000000000000000010111011000000011000101000000000010110010000000100000000000000000111000000000001000000000000000000110001010100000000000000000000") port map( O =>C_3_S_2_L_4_out, I0 =>  inp_feat(9), I1 =>  inp_feat(407), I2 =>  inp_feat(193), I3 =>  inp_feat(449), I4 =>  inp_feat(352), I5 =>  inp_feat(354), I6 =>  inp_feat(201), I7 =>  inp_feat(331)); 
C_3_S_2_L_5_inst : LUT8 generic map(INIT => "0010001000001000001000100000100000100000000010000010101010000000010000101000000000000000000000000000000000000000000000000000000010001000000000001011101100000000000010000000000000100010000010000000000000000000001000100000000000000010000000000000000010000000") port map( O =>C_3_S_2_L_5_out, I0 =>  inp_feat(452), I1 =>  inp_feat(465), I2 =>  inp_feat(362), I3 =>  inp_feat(50), I4 =>  inp_feat(463), I5 =>  inp_feat(232), I6 =>  inp_feat(298), I7 =>  inp_feat(475)); 
C_3_S_2_L_6_inst : LUT8 generic map(INIT => "1111010001110111000000010001000011010101100000001000000010000000100000100011000100000001000000000010000010000000001001101000000000000000000000000001000000000000000000001000000010000000000000001000000000000000100000001000000000000000000000000000000000000000") port map( O =>C_3_S_2_L_6_out, I0 =>  inp_feat(462), I1 =>  inp_feat(98), I2 =>  inp_feat(478), I3 =>  inp_feat(368), I4 =>  inp_feat(161), I5 =>  inp_feat(206), I6 =>  inp_feat(290), I7 =>  inp_feat(41)); 
C_3_S_2_L_7_inst : LUT8 generic map(INIT => "1010000010101011011000001000000010000000100000000000000000000000100000000100111100000000010000000000000010000000100000001100100000000010000000100000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_2_L_7_out, I0 =>  inp_feat(259), I1 =>  inp_feat(354), I2 =>  inp_feat(11), I3 =>  inp_feat(177), I4 =>  inp_feat(321), I5 =>  inp_feat(387), I6 =>  inp_feat(71), I7 =>  inp_feat(327)); 
C_3_S_3_L_0_inst : LUT8 generic map(INIT => "1001101000000000000000000000000000001010000011000000000000000000100010000000010010000000000000001000101010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010000010000000000000000000") port map( O =>C_3_S_3_L_0_out, I0 =>  inp_feat(212), I1 =>  inp_feat(458), I2 =>  inp_feat(347), I3 =>  inp_feat(110), I4 =>  inp_feat(403), I5 =>  inp_feat(258), I6 =>  inp_feat(508), I7 =>  inp_feat(311)); 
C_3_S_3_L_1_inst : LUT8 generic map(INIT => "0000000100000100000000000000000010000000000000000000000000000000000010001000000001000000000000001000100001001100000000000000000000001000000000011010010010000001000110000000010000001010010000010000001000010001000000000000010000001111010011010101111100001100") port map( O =>C_3_S_3_L_1_out, I0 =>  inp_feat(427), I1 =>  inp_feat(259), I2 =>  inp_feat(462), I3 =>  inp_feat(237), I4 =>  inp_feat(468), I5 =>  inp_feat(70), I6 =>  inp_feat(192), I7 =>  inp_feat(504)); 
C_3_S_3_L_2_inst : LUT8 generic map(INIT => "0000101000000000100010100000000000000000000000000000000000000000111110100000000000000000000000000000000000000000000000000000000010101011000000000000000000000000000000000000000000000000000000001000001100000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_3_L_2_out, I0 =>  inp_feat(376), I1 =>  inp_feat(23), I2 =>  inp_feat(508), I3 =>  inp_feat(311), I4 =>  inp_feat(191), I5 =>  inp_feat(266), I6 =>  inp_feat(478), I7 =>  inp_feat(65)); 
C_3_S_3_L_3_inst : LUT8 generic map(INIT => "1000110000101100010111000000000011001100000010000010110000001000100000000000000000000100000001000000000000001000000010001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_3_L_3_out, I0 =>  inp_feat(382), I1 =>  inp_feat(183), I2 =>  inp_feat(82), I3 =>  inp_feat(456), I4 =>  inp_feat(21), I5 =>  inp_feat(65), I6 =>  inp_feat(492), I7 =>  inp_feat(266)); 
C_3_S_3_L_4_inst : LUT8 generic map(INIT => "0010100010000000010000001011010100000000000000000000110000000000000101100000000001110000111100000000100100000001000000000100111100000000000000000000000010100000000000000000000000000000000000010000000000110000000100000001000110100000000000000000000011001111") port map( O =>C_3_S_3_L_4_out, I0 =>  inp_feat(120), I1 =>  inp_feat(275), I2 =>  inp_feat(394), I3 =>  inp_feat(126), I4 =>  inp_feat(388), I5 =>  inp_feat(5), I6 =>  inp_feat(53), I7 =>  inp_feat(77)); 
C_3_S_3_L_5_inst : LUT8 generic map(INIT => "1101000010000000011101010000001110000000000000000001011100101001111100000100000000010000000100000000000000000000000000000000000000010010000100000001000100000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_3_L_5_out, I0 =>  inp_feat(336), I1 =>  inp_feat(29), I2 =>  inp_feat(340), I3 =>  inp_feat(364), I4 =>  inp_feat(204), I5 =>  inp_feat(178), I6 =>  inp_feat(388), I7 =>  inp_feat(310)); 
C_3_S_3_L_6_inst : LUT8 generic map(INIT => "1110000011111000110100001011100000000000101100000110000011100000101010001001100011010000111010000000000001010000010000011111001000000000010000000000000000000000000000000000000001000000100010000000000000001000000000000000100000000000010010000000000010000000") port map( O =>C_3_S_3_L_6_out, I0 =>  inp_feat(451), I1 =>  inp_feat(52), I2 =>  inp_feat(148), I3 =>  inp_feat(6), I4 =>  inp_feat(247), I5 =>  inp_feat(220), I6 =>  inp_feat(83), I7 =>  inp_feat(328)); 
C_3_S_3_L_7_inst : LUT8 generic map(INIT => "1100001000100000100000100000000010101010000000001000100000001100101010100010110010101110000000000001001000000010000000110000000010010000000000000000000000000000000000000000000000000111000000001000101001000110000000000000000000001010001111000000111101001000") port map( O =>C_3_S_3_L_7_out, I0 =>  inp_feat(221), I1 =>  inp_feat(413), I2 =>  inp_feat(485), I3 =>  inp_feat(340), I4 =>  inp_feat(385), I5 =>  inp_feat(354), I6 =>  inp_feat(152), I7 =>  inp_feat(74)); 
C_3_S_4_L_0_inst : LUT8 generic map(INIT => "1000000000000010010101000000000011101000101000100101000000100000110000000100010000000000110000001100000000000000000000000000000000000000000000000000000000000000000000001010001000010000100000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_3_S_4_L_0_out, I0 =>  inp_feat(508), I1 =>  inp_feat(290), I2 =>  inp_feat(387), I3 =>  inp_feat(376), I4 =>  inp_feat(264), I5 =>  inp_feat(347), I6 =>  inp_feat(65), I7 =>  inp_feat(492)); 
C_3_S_4_L_1_inst : LUT8 generic map(INIT => "0100000100000000011101100000011000000100100000001100000000000010000000000000000000000000000000000000000000000000000000000000000000101000000000000110000000100000101010001001001011000000111100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_4_L_1_out, I0 =>  inp_feat(7), I1 =>  inp_feat(376), I2 =>  inp_feat(5), I3 =>  inp_feat(424), I4 =>  inp_feat(388), I5 =>  inp_feat(100), I6 =>  inp_feat(266), I7 =>  inp_feat(149)); 
C_3_S_4_L_2_inst : LUT8 generic map(INIT => "1110101010101010110001000000000011101000000000000000010000110000000010000000000010001000000000000000100000000000000010000011000000110001001000000101111101010000000000000000000001000001011001000100000000000000000001000111010100000000000000000100000000000000") port map( O =>C_3_S_4_L_2_out, I0 =>  inp_feat(192), I1 =>  inp_feat(259), I2 =>  inp_feat(477), I3 =>  inp_feat(178), I4 =>  inp_feat(70), I5 =>  inp_feat(478), I6 =>  inp_feat(93), I7 =>  inp_feat(253)); 
C_3_S_4_L_3_inst : LUT8 generic map(INIT => "0101000011000101010000000100010111000000011100000000000000000000000001000000000000000000110100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_4_L_3_out, I0 =>  inp_feat(473), I1 =>  inp_feat(15), I2 =>  inp_feat(321), I3 =>  inp_feat(25), I4 =>  inp_feat(390), I5 =>  inp_feat(72), I6 =>  inp_feat(157), I7 =>  inp_feat(143)); 
C_3_S_4_L_4_inst : LUT8 generic map(INIT => "0101100011010101110000000100010111000000011100000000000000000000000001000000000000000000110100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_4_L_4_out, I0 =>  inp_feat(473), I1 =>  inp_feat(15), I2 =>  inp_feat(321), I3 =>  inp_feat(25), I4 =>  inp_feat(390), I5 =>  inp_feat(72), I6 =>  inp_feat(157), I7 =>  inp_feat(143)); 
C_3_S_4_L_5_inst : LUT8 generic map(INIT => "1010000010001000100010100000000001110111000000000111001100000100000000000000000000000000000000000000000000000000001000000000000000011000100000000010001010000000000100000100000001000100010000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_3_S_4_L_5_out, I0 =>  inp_feat(209), I1 =>  inp_feat(435), I2 =>  inp_feat(337), I3 =>  inp_feat(95), I4 =>  inp_feat(53), I5 =>  inp_feat(70), I6 =>  inp_feat(143), I7 =>  inp_feat(71)); 
C_3_S_4_L_6_inst : LUT8 generic map(INIT => "0011010000000000001000001000000000000000000000000000000010000000000110010000000010000001000000000000000000000000000000000000000000000001000000000010000011000000000000000000000000000000100000000110000000000000000000000000000000000000000000000000000010000000") port map( O =>C_3_S_4_L_6_out, I0 =>  inp_feat(477), I1 =>  inp_feat(463), I2 =>  inp_feat(325), I3 =>  inp_feat(58), I4 =>  inp_feat(29), I5 =>  inp_feat(301), I6 =>  inp_feat(310), I7 =>  inp_feat(74)); 
C_3_S_4_L_7_inst : LUT8 generic map(INIT => "0001000111000000000010010010000011110100101101101011111111000001000000100010000010100000000000001100000000000000111111110000100010000000000000010000000000000000000001000000000001000101000001100000000000000000000000000000000001000000000000001001000100000000") port map( O =>C_3_S_4_L_7_out, I0 =>  inp_feat(6), I1 =>  inp_feat(420), I2 =>  inp_feat(83), I3 =>  inp_feat(373), I4 =>  inp_feat(42), I5 =>  inp_feat(82), I6 =>  inp_feat(21), I7 =>  inp_feat(327)); 
C_4_S_0_L_0_inst : LUT8 generic map(INIT => "0000000010000000000000001000000000000000000000000000000000000000100000001000000000000000100000001000000010000000000000000000000000000010000000100000000010000000101100100010000000000000000000000000000010000000000000000000000010100000100000000000000000000000") port map( O =>C_4_S_0_L_0_out, I0 =>  inp_feat(201), I1 =>  inp_feat(480), I2 =>  inp_feat(222), I3 =>  inp_feat(152), I4 =>  inp_feat(259), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_4_S_0_L_1_inst : LUT8 generic map(INIT => "1000111000000000000000000000000000000000000000000000000000000000101010100000000000001000000000000000111000000000000000000000000011010100101100000000000000000000000010100100000000000000000000001010001000000000000000000000000000001111000000000000000000000000") port map( O =>C_4_S_0_L_1_out, I0 =>  inp_feat(353), I1 =>  inp_feat(149), I2 =>  inp_feat(376), I3 =>  inp_feat(403), I4 =>  inp_feat(143), I5 =>  inp_feat(277), I6 =>  inp_feat(70), I7 =>  inp_feat(440)); 
C_4_S_0_L_2_inst : LUT8 generic map(INIT => "0001000000001000010000001000000000000000000000000000000000000000000000000000000010000000000000000010001000000000000000000001000000000000001100011001000011110011001000000011000010100001011101110010000000000000000000001100000000100000001000000000000011100000") port map( O =>C_4_S_0_L_2_out, I0 =>  inp_feat(77), I1 =>  inp_feat(158), I2 =>  inp_feat(93), I3 =>  inp_feat(70), I4 =>  inp_feat(462), I5 =>  inp_feat(83), I6 =>  inp_feat(91), I7 =>  inp_feat(65)); 
C_4_S_0_L_3_inst : LUT8 generic map(INIT => "1110100000110011001100000000000000111010000101011000100000000000110010001000000010000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_0_L_3_out, I0 =>  inp_feat(465), I1 =>  inp_feat(57), I2 =>  inp_feat(154), I3 =>  inp_feat(15), I4 =>  inp_feat(212), I5 =>  inp_feat(494), I6 =>  inp_feat(116), I7 =>  inp_feat(266)); 
C_4_S_0_L_4_inst : LUT8 generic map(INIT => "0000001000000010010010100000000010000000000010001000100000000000000000000000000000000000000000000000000000000000100000000000000010100000000000001000000000000000100000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_0_L_4_out, I0 =>  inp_feat(86), I1 =>  inp_feat(493), I2 =>  inp_feat(430), I3 =>  inp_feat(296), I4 =>  inp_feat(388), I5 =>  inp_feat(80), I6 =>  inp_feat(266), I7 =>  inp_feat(508)); 
C_4_S_0_L_5_inst : LUT8 generic map(INIT => "1101100011100000110010000000000011011111110000000100010100000000100000000000100000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000110000101000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_0_L_5_out, I0 =>  inp_feat(470), I1 =>  inp_feat(340), I2 =>  inp_feat(221), I3 =>  inp_feat(95), I4 =>  inp_feat(144), I5 =>  inp_feat(204), I6 =>  inp_feat(183), I7 =>  inp_feat(328)); 
C_4_S_0_L_6_inst : LUT8 generic map(INIT => "1001100000001010000001000000001000000000000000000000000010000000100100000001101000010010001000100000000000000000000000000000000011111000100011100100011000000010000000000000000000000000000000000100000010001010000000001010001000000000000000000000000000000000") port map( O =>C_4_S_0_L_6_out, I0 =>  inp_feat(483), I1 =>  inp_feat(31), I2 =>  inp_feat(192), I3 =>  inp_feat(70), I4 =>  inp_feat(469), I5 =>  inp_feat(143), I6 =>  inp_feat(416), I7 =>  inp_feat(275)); 
C_4_S_0_L_7_inst : LUT8 generic map(INIT => "1010000000100000011111110000000000000000101110001000100000000000110001100000000000111000000000000010000000100000000000000000000000000000000000000010001000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_0_L_7_out, I0 =>  inp_feat(52), I1 =>  inp_feat(316), I2 =>  inp_feat(5), I3 =>  inp_feat(86), I4 =>  inp_feat(442), I5 =>  inp_feat(415), I6 =>  inp_feat(310), I7 =>  inp_feat(327)); 
C_4_S_1_L_0_inst : LUT8 generic map(INIT => "0000110011101111000001100110101100000000000000000000000010000000100010001000100010000000100000000000000000000000000000000000000000001100101010101010100011110010000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_1_L_0_out, I0 =>  inp_feat(478), I1 =>  inp_feat(277), I2 =>  inp_feat(275), I3 =>  inp_feat(70), I4 =>  inp_feat(468), I5 =>  inp_feat(143), I6 =>  inp_feat(503), I7 =>  inp_feat(375)); 
C_4_S_1_L_1_inst : LUT8 generic map(INIT => "1010000000001000100000000000000001110000100000000010000000000000110000000000000010000000000000001111000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010001000000000") port map( O =>C_4_S_1_L_1_out, I0 =>  inp_feat(280), I1 =>  inp_feat(11), I2 =>  inp_feat(374), I3 =>  inp_feat(478), I4 =>  inp_feat(152), I5 =>  inp_feat(480), I6 =>  inp_feat(59), I7 =>  inp_feat(329)); 
C_4_S_1_L_2_inst : LUT8 generic map(INIT => "0010000010110000000000001110000011000000000000000000001000000000000000000000000001000000000000000101000000000000000000000000000010000000110000000000000000000000110010100000100000000000100000000000000000000000000000000000000010000000000000000000000010000000") port map( O =>C_4_S_1_L_2_out, I0 =>  inp_feat(391), I1 =>  inp_feat(386), I2 =>  inp_feat(403), I3 =>  inp_feat(376), I4 =>  inp_feat(267), I5 =>  inp_feat(508), I6 =>  inp_feat(93), I7 =>  inp_feat(65)); 
C_4_S_1_L_3_inst : LUT8 generic map(INIT => "1111000100000001010010010000000111000101100000110000000101010111000000000000000000000000000000000000000000000000000001000000000000000001000000010000000000000001000000001000000100000001000101110000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_1_L_3_out, I0 =>  inp_feat(462), I1 =>  inp_feat(388), I2 =>  inp_feat(70), I3 =>  inp_feat(95), I4 =>  inp_feat(77), I5 =>  inp_feat(158), I6 =>  inp_feat(143), I7 =>  inp_feat(93)); 
C_4_S_1_L_4_inst : LUT8 generic map(INIT => "1000100010000000110110000001000000110000000000000000100001000000100010000000000011010000010100001000000000000000000000000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000") port map( O =>C_4_S_1_L_4_out, I0 =>  inp_feat(166), I1 =>  inp_feat(201), I2 =>  inp_feat(427), I3 =>  inp_feat(41), I4 =>  inp_feat(302), I5 =>  inp_feat(414), I6 =>  inp_feat(42), I7 =>  inp_feat(327)); 
C_4_S_1_L_5_inst : LUT8 generic map(INIT => "1001010000100000000001000000000001000000000000001100000000000000000000000000000000001001000000001111100010000000110000001000000010000000000000000000000100000000010100000000000001000000001100001100010000000000000010110000000011110000000100000101000000110000") port map( O =>C_4_S_1_L_5_out, I0 =>  inp_feat(382), I1 =>  inp_feat(11), I2 =>  inp_feat(376), I3 =>  inp_feat(327), I4 =>  inp_feat(21), I5 =>  inp_feat(82), I6 =>  inp_feat(295), I7 =>  inp_feat(504)); 
C_4_S_1_L_6_inst : LUT8 generic map(INIT => "0010001100000000000000001000000000100000000000000000000000000000000000000000000010000000100010000000000000000000000000000000000000000011100000000010000100000000000000000010000000000001000000100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_1_L_6_out, I0 =>  inp_feat(445), I1 =>  inp_feat(285), I2 =>  inp_feat(511), I3 =>  inp_feat(295), I4 =>  inp_feat(392), I5 =>  inp_feat(297), I6 =>  inp_feat(403), I7 =>  inp_feat(163)); 
C_4_S_1_L_7_inst : LUT8 generic map(INIT => "1000000011000000110000000001000011000000100000000000000000000001000101101111000001110000111100010000000001000000010000001001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000") port map( O =>C_4_S_1_L_7_out, I0 =>  inp_feat(275), I1 =>  inp_feat(77), I2 =>  inp_feat(18), I3 =>  inp_feat(388), I4 =>  inp_feat(53), I5 =>  inp_feat(93), I6 =>  inp_feat(70), I7 =>  inp_feat(266)); 
C_4_S_2_L_0_inst : LUT8 generic map(INIT => "1010001000000000001000100000000011001000110000000000000000100000000000000000000000000000000100001101000010000000000000001001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_2_L_0_out, I0 =>  inp_feat(355), I1 =>  inp_feat(372), I2 =>  inp_feat(183), I3 =>  inp_feat(443), I4 =>  inp_feat(424), I5 =>  inp_feat(23), I6 =>  inp_feat(298), I7 =>  inp_feat(41)); 
C_4_S_2_L_1_inst : LUT8 generic map(INIT => "0001000000000000000000001100000000010000000000000000000000000000000010001010000000000000010001000000100000000000000000000000010001100000110000000100000000100101000000000000000100000000000000000000000011100110010101010110011110001000001101010000000001010101") port map( O =>C_4_S_2_L_1_out, I0 =>  inp_feat(158), I1 =>  inp_feat(393), I2 =>  inp_feat(468), I3 =>  inp_feat(462), I4 =>  inp_feat(427), I5 =>  inp_feat(93), I6 =>  inp_feat(388), I7 =>  inp_feat(70)); 
C_4_S_2_L_2_inst : LUT8 generic map(INIT => "0110111011100000000000000000000011100000111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_2_L_2_out, I0 =>  inp_feat(212), I1 =>  inp_feat(465), I2 =>  inp_feat(224), I3 =>  inp_feat(172), I4 =>  inp_feat(311), I5 =>  inp_feat(470), I6 =>  inp_feat(266), I7 =>  inp_feat(143)); 
C_4_S_2_L_3_inst : LUT8 generic map(INIT => "0010110100000010000011110000010000000000000000000000000000000000100010000000000000001110000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000") port map( O =>C_4_S_2_L_3_out, I0 =>  inp_feat(464), I1 =>  inp_feat(52), I2 =>  inp_feat(369), I3 =>  inp_feat(368), I4 =>  inp_feat(172), I5 =>  inp_feat(311), I6 =>  inp_feat(470), I7 =>  inp_feat(143)); 
C_4_S_2_L_4_inst : LUT8 generic map(INIT => "1011101100001010100000001001000000011010000000001100000000000000010011000000000011001111000000101110100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_4_S_2_L_4_out, I0 =>  inp_feat(149), I1 =>  inp_feat(477), I2 =>  inp_feat(201), I3 =>  inp_feat(93), I4 =>  inp_feat(70), I5 =>  inp_feat(152), I6 =>  inp_feat(480), I7 =>  inp_feat(143)); 
C_4_S_2_L_5_inst : LUT8 generic map(INIT => "0000101001000000110011110000001000000000000000000000000000000000100000000000000010001011000000000000000000000010000000010000000000100100000000110000000001001111100000000000001000000001010000010000000000000000000011010000000000000011000001100010101100000111") port map( O =>C_4_S_2_L_5_out, I0 =>  inp_feat(77), I1 =>  inp_feat(416), I2 =>  inp_feat(70), I3 =>  inp_feat(95), I4 =>  inp_feat(192), I5 =>  inp_feat(5), I6 =>  inp_feat(168), I7 =>  inp_feat(53)); 
C_4_S_2_L_6_inst : LUT8 generic map(INIT => "0110000100001111000000001000000111011010101000100000000010000000101000100010101000000000000000001110011000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_2_L_6_out, I0 =>  inp_feat(478), I1 =>  inp_feat(192), I2 =>  inp_feat(436), I3 =>  inp_feat(83), I4 =>  inp_feat(148), I5 =>  inp_feat(336), I6 =>  inp_feat(149), I7 =>  inp_feat(266)); 
C_4_S_2_L_7_inst : LUT8 generic map(INIT => "0110000010000000000100001000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000000000101000011100000000000000000000001000001101000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_2_L_7_out, I0 =>  inp_feat(5), I1 =>  inp_feat(71), I2 =>  inp_feat(298), I3 =>  inp_feat(63), I4 =>  inp_feat(310), I5 =>  inp_feat(74), I6 =>  inp_feat(91), I7 =>  inp_feat(149)); 
C_4_S_3_L_0_inst : LUT8 generic map(INIT => "1001100000000100100010000010000000000000000000001100111000000000100010001000000010001000001000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_3_L_0_out, I0 =>  inp_feat(424), I1 =>  inp_feat(376), I2 =>  inp_feat(443), I3 =>  inp_feat(297), I4 =>  inp_feat(181), I5 =>  inp_feat(116), I6 =>  inp_feat(83), I7 =>  inp_feat(143)); 
C_4_S_3_L_1_inst : LUT8 generic map(INIT => "1100001000001010001110000100100011110000001000010000010000001000000000000000000000000000000000000000000000100010000000000000000010000000000000000000000000000000101000000000000000000000000100000000000000000000000000000000000001001000000000000000000000000010") port map( O =>C_4_S_3_L_1_out, I0 =>  inp_feat(427), I1 =>  inp_feat(11), I2 =>  inp_feat(441), I3 =>  inp_feat(212), I4 =>  inp_feat(381), I5 =>  inp_feat(268), I6 =>  inp_feat(311), I7 =>  inp_feat(290)); 
C_4_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000011000100000000010000000000000000000100000010000010000000000000000000000001001101000000000000000000000010000000000000000000000000100100000000000000000000000000001111111101100111110010000101001100000100000011100000000000000000") port map( O =>C_4_S_3_L_2_out, I0 =>  inp_feat(362), I1 =>  inp_feat(499), I2 =>  inp_feat(25), I3 =>  inp_feat(156), I4 =>  inp_feat(250), I5 =>  inp_feat(455), I6 =>  inp_feat(465), I7 =>  inp_feat(122)); 
C_4_S_3_L_3_inst : LUT8 generic map(INIT => "0101110100000000111111000000000000000000000000000100000000000000110011000000000001001000000010001000000000001100010110000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_3_L_3_out, I0 =>  inp_feat(318), I1 =>  inp_feat(212), I2 =>  inp_feat(170), I3 =>  inp_feat(349), I4 =>  inp_feat(6), I5 =>  inp_feat(148), I6 =>  inp_feat(83), I7 =>  inp_feat(143)); 
C_4_S_3_L_4_inst : LUT8 generic map(INIT => "1000110101001001000000000000000000000000010000110000000000001000101111010010101000010000001000000000010000000000000000000000000000101100001000000000000000000010000000000000000000000000000000000110100010001011000010000010001000000000001000010000000010000011") port map( O =>C_4_S_3_L_4_out, I0 =>  inp_feat(201), I1 =>  inp_feat(367), I2 =>  inp_feat(295), I3 =>  inp_feat(6), I4 =>  inp_feat(415), I5 =>  inp_feat(148), I6 =>  inp_feat(331), I7 =>  inp_feat(161)); 
C_4_S_3_L_5_inst : LUT8 generic map(INIT => "0000000001001111001000000101011000000100010000000000001001000000000010100000110001010010010001000000001000001010000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000") port map( O =>C_4_S_3_L_5_out, I0 =>  inp_feat(100), I1 =>  inp_feat(382), I2 =>  inp_feat(42), I3 =>  inp_feat(65), I4 =>  inp_feat(149), I5 =>  inp_feat(35), I6 =>  inp_feat(507), I7 =>  inp_feat(266)); 
C_4_S_3_L_6_inst : LUT8 generic map(INIT => "1000110001001000000000000000000000000000000000000000001010000000110000000010000010000000000000000000000010000000000010110000000100001000000000000000000010000000000001000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000") port map( O =>C_4_S_3_L_6_out, I0 =>  inp_feat(259), I1 =>  inp_feat(203), I2 =>  inp_feat(201), I3 =>  inp_feat(100), I4 =>  inp_feat(267), I5 =>  inp_feat(21), I6 =>  inp_feat(65), I7 =>  inp_feat(328)); 
C_4_S_3_L_7_inst : LUT8 generic map(INIT => "0110101110010000010001100000000011000000000110010000000000000000000000001100000000000100000000000000001110000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_3_L_7_out, I0 =>  inp_feat(120), I1 =>  inp_feat(388), I2 =>  inp_feat(510), I3 =>  inp_feat(408), I4 =>  inp_feat(144), I5 =>  inp_feat(297), I6 =>  inp_feat(392), I7 =>  inp_feat(403)); 
C_4_S_4_L_0_inst : LUT8 generic map(INIT => "1100011000000011001011111000001000000000010010000000011000111011000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_4_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(91), I2 =>  inp_feat(82), I3 =>  inp_feat(507), I4 =>  inp_feat(65), I5 =>  inp_feat(415), I6 =>  inp_feat(266), I7 =>  inp_feat(143)); 
C_4_S_4_L_1_inst : LUT8 generic map(INIT => "0010000000010000000000000000000101010000111101110100000011110011000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_4_L_1_out, I0 =>  inp_feat(192), I1 =>  inp_feat(342), I2 =>  inp_feat(393), I3 =>  inp_feat(126), I4 =>  inp_feat(125), I5 =>  inp_feat(70), I6 =>  inp_feat(266), I7 =>  inp_feat(143)); 
C_4_S_4_L_2_inst : LUT8 generic map(INIT => "1011001010101010011111111010100010100000000001000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_4_L_2_out, I0 =>  inp_feat(201), I1 =>  inp_feat(6), I2 =>  inp_feat(480), I3 =>  inp_feat(70), I4 =>  inp_feat(152), I5 =>  inp_feat(310), I6 =>  inp_feat(266), I7 =>  inp_feat(143)); 
C_4_S_4_L_3_inst : LUT8 generic map(INIT => "0100010100001010010000000000000011010100000010000000000000000000000000000000000000000000000000000000001000000000000000000000000011011100001010101000000000000000110001000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000") port map( O =>C_4_S_4_L_3_out, I0 =>  inp_feat(70), I1 =>  inp_feat(480), I2 =>  inp_feat(375), I3 =>  inp_feat(108), I4 =>  inp_feat(328), I5 =>  inp_feat(273), I6 =>  inp_feat(169), I7 =>  inp_feat(347)); 
C_4_S_4_L_4_inst : LUT8 generic map(INIT => "1110101000000000101010000010000001110000000000000011000000000000000110110001000110100111001000000000000000000000000000000000001001000001000000000010000010000000000000000000000000111010000000000100010000000010101010000010001100000001000000000010111100100000") port map( O =>C_4_S_4_L_4_out, I0 =>  inp_feat(420), I1 =>  inp_feat(206), I2 =>  inp_feat(162), I3 =>  inp_feat(327), I4 =>  inp_feat(74), I5 =>  inp_feat(480), I6 =>  inp_feat(367), I7 =>  inp_feat(52)); 
C_4_S_4_L_5_inst : LUT8 generic map(INIT => "1010000000000000000100000110000011011000000010001111100111110000000000000000000000000000000000000000000000000000000000000000000001000010000000000010000000000000000000000000000011001011000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_4_L_5_out, I0 =>  inp_feat(290), I1 =>  inp_feat(11), I2 =>  inp_feat(447), I3 =>  inp_feat(68), I4 =>  inp_feat(385), I5 =>  inp_feat(508), I6 =>  inp_feat(266), I7 =>  inp_feat(141)); 
C_4_S_4_L_6_inst : LUT8 generic map(INIT => "1000010110011000001000000000000000000000010000001000000010000000000001110100010000100000000000010000010000000000000000001000000000000000000010000000010010000000000001100000000000000000100000000000000000000001000000011000000100000001000000000000000000000000") port map( O =>C_4_S_4_L_6_out, I0 =>  inp_feat(302), I1 =>  inp_feat(154), I2 =>  inp_feat(318), I3 =>  inp_feat(344), I4 =>  inp_feat(303), I5 =>  inp_feat(1), I6 =>  inp_feat(238), I7 =>  inp_feat(448)); 
C_4_S_4_L_7_inst : LUT8 generic map(INIT => "1010010010001100000000000000010001100000100000000000000000000000100001000010010000000000000000000000000000000000000000000000000010001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_4_S_4_L_7_out, I0 =>  inp_feat(191), I1 =>  inp_feat(368), I2 =>  inp_feat(198), I3 =>  inp_feat(508), I4 =>  inp_feat(311), I5 =>  inp_feat(116), I6 =>  inp_feat(471), I7 =>  inp_feat(71)); 
C_5_S_0_L_0_inst : LUT8 generic map(INIT => "0000001000000010001000000010000000000000000000000000000000000000101000100000000000000000000010100000000000000000000000100000001000001000000010000000100000000010000000000000000000000000000000000010101000000000100000000000000000000000000000000000000000000000") port map( O =>C_5_S_0_L_0_out, I0 =>  inp_feat(10), I1 =>  inp_feat(462), I2 =>  inp_feat(158), I3 =>  inp_feat(427), I4 =>  inp_feat(224), I5 =>  inp_feat(30), I6 =>  inp_feat(70), I7 =>  inp_feat(503)); 
C_5_S_0_L_1_inst : LUT8 generic map(INIT => "1110010011001000111000001100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000001010000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000") port map( O =>C_5_S_0_L_1_out, I0 =>  inp_feat(443), I1 =>  inp_feat(386), I2 =>  inp_feat(277), I3 =>  inp_feat(21), I4 =>  inp_feat(17), I5 =>  inp_feat(242), I6 =>  inp_feat(214), I7 =>  inp_feat(15)); 
C_5_S_0_L_2_inst : LUT8 generic map(INIT => "1000000110000000000000001010101010000000110000000000000000100000000001000010000000000000001000000001000000000000000000000000000010100010100000000000000000000000000000001100000000000000000000000000000000000000000000000000000010100000000000000000000000000000") port map( O =>C_5_S_0_L_2_out, I0 =>  inp_feat(340), I1 =>  inp_feat(87), I2 =>  inp_feat(328), I3 =>  inp_feat(465), I4 =>  inp_feat(15), I5 =>  inp_feat(77), I6 =>  inp_feat(387), I7 =>  inp_feat(70)); 
C_5_S_0_L_3_inst : LUT8 generic map(INIT => "1101001100001111111101010000010100000001000011110000010000000101110100100000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000010000000100000001") port map( O =>C_5_S_0_L_3_out, I0 =>  inp_feat(29), I1 =>  inp_feat(6), I2 =>  inp_feat(442), I3 =>  inp_feat(340), I4 =>  inp_feat(65), I5 =>  inp_feat(251), I6 =>  inp_feat(492), I7 =>  inp_feat(327)); 
C_5_S_0_L_4_inst : LUT8 generic map(INIT => "0000000001001000000010000000000000101000000000001000001010000000100010101100111000001000010010001100110011101110100010001100100010011000000000000000001000000000000000000000000010001000100010000000000000001000000000000000000000000000000000001000100010001000") port map( O =>C_5_S_0_L_4_out, I0 =>  inp_feat(41), I1 =>  inp_feat(201), I2 =>  inp_feat(420), I3 =>  inp_feat(475), I4 =>  inp_feat(65), I5 =>  inp_feat(498), I6 =>  inp_feat(152), I7 =>  inp_feat(168)); 
C_5_S_0_L_5_inst : LUT8 generic map(INIT => "1000110011001100100000001000000000000000000000000000000000000000100010000001000000100000000000001000000000000000000000000000000011010000000110001000101000000000000000000000000000000000000000001101000001010000001110110000101010000000000000000000000000000000") port map( O =>C_5_S_0_L_5_out, I0 =>  inp_feat(478), I1 =>  inp_feat(93), I2 =>  inp_feat(365), I3 =>  inp_feat(373), I4 =>  inp_feat(178), I5 =>  inp_feat(8), I6 =>  inp_feat(100), I7 =>  inp_feat(34)); 
C_5_S_0_L_6_inst : LUT8 generic map(INIT => "1010100000001000101000000000000010000000100000001010000001000000000000001000001010001000100010000100100010000010100010001100101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000001000") port map( O =>C_5_S_0_L_6_out, I0 =>  inp_feat(43), I1 =>  inp_feat(384), I2 =>  inp_feat(115), I3 =>  inp_feat(433), I4 =>  inp_feat(151), I5 =>  inp_feat(362), I6 =>  inp_feat(3), I7 =>  inp_feat(188)); 
C_5_S_0_L_7_inst : LUT8 generic map(INIT => "1110101100001000001010000000000000000001000000000000000010110000000000111000001000001100000000000000000000000000000000000000000010000010000000001010101110101010000000000000010001010100010001000001101100000000000001110000000000000000000000000000000101000000") port map( O =>C_5_S_0_L_7_out, I0 =>  inp_feat(289), I1 =>  inp_feat(295), I2 =>  inp_feat(382), I3 =>  inp_feat(181), I4 =>  inp_feat(65), I5 =>  inp_feat(116), I6 =>  inp_feat(494), I7 =>  inp_feat(498)); 
C_5_S_1_L_0_inst : LUT8 generic map(INIT => "1010000010101000101010001000000010000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000001010000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_5_S_1_L_0_out, I0 =>  inp_feat(54), I1 =>  inp_feat(264), I2 =>  inp_feat(183), I3 =>  inp_feat(27), I4 =>  inp_feat(173), I5 =>  inp_feat(387), I6 =>  inp_feat(214), I7 =>  inp_feat(15)); 
C_5_S_1_L_1_inst : LUT8 generic map(INIT => "0010100000011000011010000000000010001010000010000000000000000000101010001100000000001000000000000000000000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000010000000000000011000000000000000000000000000000000000000000") port map( O =>C_5_S_1_L_1_out, I0 =>  inp_feat(11), I1 =>  inp_feat(328), I2 =>  inp_feat(465), I3 =>  inp_feat(387), I4 =>  inp_feat(396), I5 =>  inp_feat(15), I6 =>  inp_feat(207), I7 =>  inp_feat(46)); 
C_5_S_1_L_2_inst : LUT8 generic map(INIT => "1010101000000000000000000000000000100000001010000011000000101000101000100000100000000000000000000000001100000000000000100000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_5_S_1_L_2_out, I0 =>  inp_feat(277), I1 =>  inp_feat(135), I2 =>  inp_feat(177), I3 =>  inp_feat(340), I4 =>  inp_feat(178), I5 =>  inp_feat(272), I6 =>  inp_feat(387), I7 =>  inp_feat(15)); 
C_5_S_1_L_3_inst : LUT8 generic map(INIT => "0100000010000000000000000100000000010000000000001100000001000000000000000000000000000000000000000000000000000000000000000100000010000000000000000100000011000000000100000000000011110000010000000000100000000000001100000000000000000000000000000001000000000000") port map( O =>C_5_S_1_L_3_out, I0 =>  inp_feat(82), I1 =>  inp_feat(394), I2 =>  inp_feat(386), I3 =>  inp_feat(432), I4 =>  inp_feat(65), I5 =>  inp_feat(295), I6 =>  inp_feat(327), I7 =>  inp_feat(83)); 
C_5_S_1_L_4_inst : LUT8 generic map(INIT => "0000001100001010000000100000000000011111100010100011111100001010101010100000000000000000000000001010111000000000000011100000100000000000000010100000100000000010000001100000000000000010000000100000000000000000000000000000100000000000000000000000111100001100") port map( O =>C_5_S_1_L_4_out, I0 =>  inp_feat(466), I1 =>  inp_feat(57), I2 =>  inp_feat(408), I3 =>  inp_feat(374), I4 =>  inp_feat(311), I5 =>  inp_feat(198), I6 =>  inp_feat(508), I7 =>  inp_feat(143)); 
C_5_S_1_L_5_inst : LUT8 generic map(INIT => "0000100011010100100000000000000000000000000000000000000000000000001000000100100000000000000000000000000000000000000000001000000001010100101110110000000000000000000000000000000000000000000000011001000011111000100000001100000000000000000001010000000100000101") port map( O =>C_5_S_1_L_5_out, I0 =>  inp_feat(6), I1 =>  inp_feat(340), I2 =>  inp_feat(120), I3 =>  inp_feat(82), I4 =>  inp_feat(181), I5 =>  inp_feat(116), I6 =>  inp_feat(65), I7 =>  inp_feat(498)); 
C_5_S_1_L_6_inst : LUT8 generic map(INIT => "0110010001000000100000000000000000000000000000000010000000000000101000010100100011100000000000001010000010100000111000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000") port map( O =>C_5_S_1_L_6_out, I0 =>  inp_feat(364), I1 =>  inp_feat(444), I2 =>  inp_feat(424), I3 =>  inp_feat(49), I4 =>  inp_feat(195), I5 =>  inp_feat(13), I6 =>  inp_feat(23), I7 =>  inp_feat(214)); 
C_5_S_1_L_7_inst : LUT8 generic map(INIT => "1110001100010110010111011001111100000000000000001000100101000001010011000101011011111111111111110000000000000000000010110000001100000001000000000000100110000111000000000000000000000000000000000000000000000000100010100000011000000000000000001000101000100011") port map( O =>C_5_S_1_L_7_out, I0 =>  inp_feat(170), I1 =>  inp_feat(212), I2 =>  inp_feat(98), I3 =>  inp_feat(100), I4 =>  inp_feat(198), I5 =>  inp_feat(466), I6 =>  inp_feat(508), I7 =>  inp_feat(124)); 
C_5_S_2_L_0_inst : LUT8 generic map(INIT => "0100010110000000000000000000000011101100000000000000000000000000110000000000000000000000000000000100110010000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000111001001100") port map( O =>C_5_S_2_L_0_out, I0 =>  inp_feat(369), I1 =>  inp_feat(354), I2 =>  inp_feat(305), I3 =>  inp_feat(452), I4 =>  inp_feat(89), I5 =>  inp_feat(465), I6 =>  inp_feat(402), I7 =>  inp_feat(15)); 
C_5_S_2_L_1_inst : LUT8 generic map(INIT => "1010100000100000001000000000000010101000101000000000000000000000111000000000000000000000000000001010000011100000000100000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000001000000010000") port map( O =>C_5_S_2_L_1_out, I0 =>  inp_feat(484), I1 =>  inp_feat(407), I2 =>  inp_feat(1), I3 =>  inp_feat(305), I4 =>  inp_feat(89), I5 =>  inp_feat(465), I6 =>  inp_feat(402), I7 =>  inp_feat(15)); 
C_5_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000100000100011000000000000000000000000000000000000000000110100000001000010101100111010000000000000000000000000000000000010100000000000001000100111101101000000000000000000000000000000001000000000000100110110011111111100000000000000000000000000000000") port map( O =>C_5_S_2_L_2_out, I0 =>  inp_feat(178), I1 =>  inp_feat(93), I2 =>  inp_feat(259), I3 =>  inp_feat(478), I4 =>  inp_feat(53), I5 =>  inp_feat(214), I6 =>  inp_feat(192), I7 =>  inp_feat(70)); 
C_5_S_2_L_3_inst : LUT8 generic map(INIT => "1101000000000000001000000000000011000000000000000100000000000000101100100000000010000010000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000") port map( O =>C_5_S_2_L_3_out, I0 =>  inp_feat(407), I1 =>  inp_feat(321), I2 =>  inp_feat(392), I3 =>  inp_feat(403), I4 =>  inp_feat(222), I5 =>  inp_feat(386), I6 =>  inp_feat(23), I7 =>  inp_feat(214)); 
C_5_S_2_L_4_inst : LUT8 generic map(INIT => "0111111000000000110000000001000011001100000000000000000000010000000000000000000000000000000000000101010101000101000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100000000000000000000") port map( O =>C_5_S_2_L_4_out, I0 =>  inp_feat(347), I1 =>  inp_feat(438), I2 =>  inp_feat(173), I3 =>  inp_feat(328), I4 =>  inp_feat(442), I5 =>  inp_feat(407), I6 =>  inp_feat(24), I7 =>  inp_feat(424)); 
C_5_S_2_L_5_inst : LUT8 generic map(INIT => "0101100110001000011000001000000001000101100000000000000000000000110010000100000010000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_5_S_2_L_5_out, I0 =>  inp_feat(27), I1 =>  inp_feat(89), I2 =>  inp_feat(290), I3 =>  inp_feat(272), I4 =>  inp_feat(298), I5 =>  inp_feat(387), I6 =>  inp_feat(508), I7 =>  inp_feat(124)); 
C_5_S_2_L_6_inst : LUT8 generic map(INIT => "0000000010010000000000000000000000000000101100010100100100000100000000000000000000000000000000000000000000000001000001000000000000011010001011111011001110101010000011011010111110111111101111110000000001000010000000000000101000010000000101011101111110001111") port map( O =>C_5_S_2_L_6_out, I0 =>  inp_feat(379), I1 =>  inp_feat(77), I2 =>  inp_feat(192), I3 =>  inp_feat(275), I4 =>  inp_feat(416), I5 =>  inp_feat(388), I6 =>  inp_feat(93), I7 =>  inp_feat(70)); 
C_5_S_2_L_7_inst : LUT8 generic map(INIT => "0010001010100011101010100000000011110011101111010000000000000000110000000110010000000000000000001010101110110011000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000") port map( O =>C_5_S_2_L_7_out, I0 =>  inp_feat(154), I1 =>  inp_feat(135), I2 =>  inp_feat(198), I3 =>  inp_feat(362), I4 =>  inp_feat(95), I5 =>  inp_feat(151), I6 =>  inp_feat(210), I7 =>  inp_feat(188)); 
C_5_S_3_L_0_inst : LUT8 generic map(INIT => "1011110110001001100000011000000111001100100111011000000110000001000000000000000000000000000000001001000000000001000000000000000000000000000000000000000100000000000000000000100000000000000000000000000001000000000000000000000000000000100000000000000000000000") port map( O =>C_5_S_3_L_0_out, I0 =>  inp_feat(272), I1 =>  inp_feat(75), I2 =>  inp_feat(336), I3 =>  inp_feat(275), I4 =>  inp_feat(354), I5 =>  inp_feat(78), I6 =>  inp_feat(452), I7 =>  inp_feat(387)); 
C_5_S_3_L_1_inst : LUT8 generic map(INIT => "1000001000000010000100000011010100000000000000100000000000000000101000011000010000100000010000000000000000000000000000000000000010000010000000000000100000110011000000000000011000000000000000001000100000000010100010001000101100000000010101000000000001000011") port map( O =>C_5_S_3_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(494), I2 =>  inp_feat(382), I3 =>  inp_feat(261), I4 =>  inp_feat(295), I5 =>  inp_feat(259), I6 =>  inp_feat(65), I7 =>  inp_feat(498)); 
C_5_S_3_L_2_inst : LUT8 generic map(INIT => "1010000000100011000001001100000010000010000000110000000000000000111111111000000010000000000001000000110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000") port map( O =>C_5_S_3_L_2_out, I0 =>  inp_feat(29), I1 =>  inp_feat(17), I2 =>  inp_feat(407), I3 =>  inp_feat(302), I4 =>  inp_feat(139), I5 =>  inp_feat(386), I6 =>  inp_feat(23), I7 =>  inp_feat(214)); 
C_5_S_3_L_3_inst : LUT8 generic map(INIT => "0100000000001000001000001000100000000000100000101011101010101010001100100000000001000000000000000000110000001100011000000000000000000100101010000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000001000000000000") port map( O =>C_5_S_3_L_3_out, I0 =>  inp_feat(340), I1 =>  inp_feat(385), I2 =>  inp_feat(21), I3 =>  inp_feat(181), I4 =>  inp_feat(79), I5 =>  inp_feat(292), I6 =>  inp_feat(374), I7 =>  inp_feat(466)); 
C_5_S_3_L_4_inst : LUT8 generic map(INIT => "1010101100000001110101000000000010010001000111110001010100110011000010000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000001000010000000000000001100110000000000000000000000000000000000000100000001010000010000000000") port map( O =>C_5_S_3_L_4_out, I0 =>  inp_feat(60), I1 =>  inp_feat(503), I2 =>  inp_feat(487), I3 =>  inp_feat(233), I4 =>  inp_feat(224), I5 =>  inp_feat(442), I6 =>  inp_feat(341), I7 =>  inp_feat(143)); 
C_5_S_3_L_5_inst : LUT8 generic map(INIT => "0110001000001000001101100000000000000000001000000000000000000000000010000000000100001111001000000000000000000000000000110000000000101011001011100010001110000010100000001000000000000010000000000011001000110101001110111111011100100010000111110000111110110111") port map( O =>C_5_S_3_L_5_out, I0 =>  inp_feat(259), I1 =>  inp_feat(192), I2 =>  inp_feat(462), I3 =>  inp_feat(416), I4 =>  inp_feat(77), I5 =>  inp_feat(93), I6 =>  inp_feat(469), I7 =>  inp_feat(70)); 
C_5_S_3_L_6_inst : LUT8 generic map(INIT => "1000100010001000010000001011100001001000000010000000000010000000000000000000000000000000000000000000100000000000000000000000000011001000110011001010000010000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000") port map( O =>C_5_S_3_L_6_out, I0 =>  inp_feat(212), I1 =>  inp_feat(397), I2 =>  inp_feat(57), I3 =>  inp_feat(268), I4 =>  inp_feat(65), I5 =>  inp_feat(407), I6 =>  inp_feat(24), I7 =>  inp_feat(292)); 
C_5_S_3_L_7_inst : LUT8 generic map(INIT => "1101100001010000100011100000110011100000000011000000110000011100000000000001000000000000000000000000000000000000001101000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001") port map( O =>C_5_S_3_L_7_out, I0 =>  inp_feat(100), I1 =>  inp_feat(383), I2 =>  inp_feat(183), I3 =>  inp_feat(479), I4 =>  inp_feat(478), I5 =>  inp_feat(176), I6 =>  inp_feat(481), I7 =>  inp_feat(188)); 
C_5_S_4_L_0_inst : LUT8 generic map(INIT => "1010000000001000000000000000010000000100000000000010000000001101000010000000000000000000000000001010110000001000000000000000000010101000000010000000000000000000000011000000010000001110000011011100110000001100000000000000000000001100000011000000000000000000") port map( O =>C_5_S_4_L_0_out, I0 =>  inp_feat(77), I1 =>  inp_feat(290), I2 =>  inp_feat(23), I3 =>  inp_feat(237), I4 =>  inp_feat(296), I5 =>  inp_feat(407), I6 =>  inp_feat(305), I7 =>  inp_feat(70)); 
C_5_S_4_L_1_inst : LUT8 generic map(INIT => "1110100100001000011010000000000001001011000000111010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000001000000000") port map( O =>C_5_S_4_L_1_out, I0 =>  inp_feat(238), I1 =>  inp_feat(494), I2 =>  inp_feat(176), I3 =>  inp_feat(464), I4 =>  inp_feat(151), I5 =>  inp_feat(210), I6 =>  inp_feat(188), I7 =>  inp_feat(288)); 
C_5_S_4_L_2_inst : LUT8 generic map(INIT => "1000000001000000010000000000000001100001110100000001000100100100110100000000010000000000000000001111111100010000101011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000") port map( O =>C_5_S_4_L_2_out, I0 =>  inp_feat(362), I1 =>  inp_feat(298), I2 =>  inp_feat(87), I3 =>  inp_feat(427), I4 =>  inp_feat(154), I5 =>  inp_feat(309), I6 =>  inp_feat(433), I7 =>  inp_feat(188)); 
C_5_S_4_L_3_inst : LUT8 generic map(INIT => "0010001010101000101000100000000000110010011000101011101010011100110000100000000000000010000000000010011000101010001010110001111000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000") port map( O =>C_5_S_4_L_3_out, I0 =>  inp_feat(179), I1 =>  inp_feat(192), I2 =>  inp_feat(401), I3 =>  inp_feat(198), I4 =>  inp_feat(362), I5 =>  inp_feat(151), I6 =>  inp_feat(210), I7 =>  inp_feat(188)); 
C_5_S_4_L_4_inst : LUT8 generic map(INIT => "1000000000000000000010000100110000000000000000000000000000000000100100000000100100010000110110000000000000000000100000001000000010001001100010011000100110001001100000000000000010000000000010000001000110010101100000011101110110000000001100010000000011010101") port map( O =>C_5_S_4_L_4_out, I0 =>  inp_feat(478), I1 =>  inp_feat(5), I2 =>  inp_feat(270), I3 =>  inp_feat(111), I4 =>  inp_feat(77), I5 =>  inp_feat(93), I6 =>  inp_feat(469), I7 =>  inp_feat(70)); 
C_5_S_4_L_5_inst : LUT8 generic map(INIT => "0010110000010001100001010000010000000000000000000101001000110000000000000000000010000000110000001010000010101000111101101010000110100001010000001000010100000000100000000100000010000000000000001000000000000000100000000000000000000000000000001000000000000000") port map( O =>C_5_S_4_L_5_out, I0 =>  inp_feat(303), I1 =>  inp_feat(373), I2 =>  inp_feat(509), I3 =>  inp_feat(87), I4 =>  inp_feat(435), I5 =>  inp_feat(507), I6 =>  inp_feat(34), I7 =>  inp_feat(83)); 
C_5_S_4_L_6_inst : LUT8 generic map(INIT => "1000011011100111100010111111111111101010001000000000000000100000101100001010000010100000101000000000000000000000000000000000000000000100000000000000000011100010000010000001000000000000000000001011000000100000001000000000000000100100000000001110010000000000") port map( O =>C_5_S_4_L_6_out, I0 =>  inp_feat(306), I1 =>  inp_feat(102), I2 =>  inp_feat(224), I3 =>  inp_feat(385), I4 =>  inp_feat(85), I5 =>  inp_feat(340), I6 =>  inp_feat(508), I7 =>  inp_feat(466)); 
C_5_S_4_L_7_inst : LUT8 generic map(INIT => "0001010000001100000000000000000001000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000010101000000010001000000000000000100110000000000000010000000000000100000000000000000000000000000000001000000000000000000000000000") port map( O =>C_5_S_4_L_7_out, I0 =>  inp_feat(371), I1 =>  inp_feat(92), I2 =>  inp_feat(484), I3 =>  inp_feat(103), I4 =>  inp_feat(116), I5 =>  inp_feat(416), I6 =>  inp_feat(424), I7 =>  inp_feat(65)); 
C_6_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_0_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_1_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_2_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_3_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_6_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_6_S_4_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(3), I3 =>  inp_feat(192), I4 =>  inp_feat(408), I5 =>  inp_feat(508), I6 =>  inp_feat(498), I7 =>  inp_feat(215)); 
C_7_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000011000000100000000000000000000000000000000000000000000000000000001101000011000000000000000000000000000000110000000000000000000000001000001100110000000000000000000100000010000000000000000000000000000000110000000000000000000000") port map( O =>C_7_S_0_L_0_out, I0 =>  inp_feat(347), I1 =>  inp_feat(466), I2 =>  inp_feat(243), I3 =>  inp_feat(462), I4 =>  inp_feat(90), I5 =>  inp_feat(508), I6 =>  inp_feat(170), I7 =>  inp_feat(215)); 
C_7_S_0_L_1_inst : LUT8 generic map(INIT => "1110001001110100011000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101010101100001010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_0_L_1_out, I0 =>  inp_feat(70), I1 =>  inp_feat(440), I2 =>  inp_feat(466), I3 =>  inp_feat(508), I4 =>  inp_feat(143), I5 =>  inp_feat(251), I6 =>  inp_feat(277), I7 =>  inp_feat(503)); 
C_7_S_0_L_2_inst : LUT8 generic map(INIT => "1000000010000000000000001000000011100000001000000011000000100000000000000010000000000000000000000000000000000000010000000101000010000000100010000010000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000001010000") port map( O =>C_7_S_0_L_2_out, I0 =>  inp_feat(308), I1 =>  inp_feat(436), I2 =>  inp_feat(15), I3 =>  inp_feat(319), I4 =>  inp_feat(480), I5 =>  inp_feat(65), I6 =>  inp_feat(221), I7 =>  inp_feat(478)); 
C_7_S_0_L_3_inst : LUT8 generic map(INIT => "0001010001001000000000000000000000111010000000100000000000000000000000000000000000000000000000000010000000000000000000000000000011011100100100000000000000000000111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_0_L_3_out, I0 =>  inp_feat(504), I1 =>  inp_feat(494), I2 =>  inp_feat(173), I3 =>  inp_feat(354), I4 =>  inp_feat(242), I5 =>  inp_feat(78), I6 =>  inp_feat(259), I7 =>  inp_feat(498)); 
C_7_S_0_L_4_inst : LUT8 generic map(INIT => "0011000000000010000001000000000011110000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000011101001011000100110001001100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_0_L_4_out, I0 =>  inp_feat(385), I1 =>  inp_feat(70), I2 =>  inp_feat(60), I3 =>  inp_feat(41), I4 =>  inp_feat(327), I5 =>  inp_feat(59), I6 =>  inp_feat(306), I7 =>  inp_feat(503)); 
C_7_S_0_L_5_inst : LUT8 generic map(INIT => "1011100010000000000010000000000010101000001000000000000000000000000000000000100000001000000000000000100010001010000000000000000010101000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_0_L_5_out, I0 =>  inp_feat(430), I1 =>  inp_feat(128), I2 =>  inp_feat(16), I3 =>  inp_feat(11), I4 =>  inp_feat(259), I5 =>  inp_feat(498), I6 =>  inp_feat(56), I7 =>  inp_feat(427)); 
C_7_S_0_L_6_inst : LUT8 generic map(INIT => "1000111010110000000000000101000100000000000000000000000000000000000011000000000000000000000000010000000000000000000000000000000010001000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_0_L_6_out, I0 =>  inp_feat(41), I1 =>  inp_feat(209), I2 =>  inp_feat(88), I3 =>  inp_feat(401), I4 =>  inp_feat(115), I5 =>  inp_feat(242), I6 =>  inp_feat(288), I7 =>  inp_feat(459)); 
C_7_S_0_L_7_inst : LUT8 generic map(INIT => "1100000000001110100000000000010110101110000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000010000000000000001000100110000000000000000000000000000001100000011000100000000001100010000000000000000000000000000000000") port map( O =>C_7_S_0_L_7_out, I0 =>  inp_feat(503), I1 =>  inp_feat(340), I2 =>  inp_feat(468), I3 =>  inp_feat(11), I4 =>  inp_feat(493), I5 =>  inp_feat(173), I6 =>  inp_feat(327), I7 =>  inp_feat(258)); 
C_7_S_1_L_0_inst : LUT8 generic map(INIT => "0101000010001000000000000000000001001000000010000100000000000000001000000000000000000000000000001100010000000000000000000000000001001000000000000000000000000000110001001000100001000000000000001100000000000000000000000000000011000100000000000000000000000000") port map( O =>C_7_S_1_L_0_out, I0 =>  inp_feat(260), I1 =>  inp_feat(86), I2 =>  inp_feat(149), I3 =>  inp_feat(478), I4 =>  inp_feat(452), I5 =>  inp_feat(508), I6 =>  inp_feat(305), I7 =>  inp_feat(215)); 
C_7_S_1_L_1_inst : LUT8 generic map(INIT => "1101000111000000110100000100000010000000000000000000000001000000100000000000000000000000010000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000") port map( O =>C_7_S_1_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(259), I2 =>  inp_feat(450), I3 =>  inp_feat(11), I4 =>  inp_feat(59), I5 =>  inp_feat(180), I6 =>  inp_feat(178), I7 =>  inp_feat(387)); 
C_7_S_1_L_2_inst : LUT8 generic map(INIT => "0111100000001000000000000000000001000000000000000000000000000000111000001000010000000000000000000000000000000000000000000000000001110000110111000000000000000000000000001000000000000000000000001111000001010000000000000000000011010000000000000000000000000000") port map( O =>C_7_S_1_L_2_out, I0 =>  inp_feat(170), I1 =>  inp_feat(258), I2 =>  inp_feat(302), I3 =>  inp_feat(475), I4 =>  inp_feat(277), I5 =>  inp_feat(212), I6 =>  inp_feat(100), I7 =>  inp_feat(440)); 
C_7_S_1_L_3_inst : LUT8 generic map(INIT => "1100010000101101110100001100000011010000000010011100000000000000000000000000000000000000000000000000000000000001000000000000000001000001010000001000000000000000110001100100001000000000000000000000000000000000000001000000000000000001000000010000000000000000") port map( O =>C_7_S_1_L_3_out, I0 =>  inp_feat(98), I1 =>  inp_feat(493), I2 =>  inp_feat(68), I3 =>  inp_feat(427), I4 =>  inp_feat(65), I5 =>  inp_feat(503), I6 =>  inp_feat(306), I7 =>  inp_feat(468)); 
C_7_S_1_L_4_inst : LUT8 generic map(INIT => "1110001011010000011100000001000011000000000000000100000001000000101000001010000000000100010100000000000000000000000000000000000000000001000000000100000000000010000000000000000000000000000000000000000000000000000000000011001000000000000000000000000000000000") port map( O =>C_7_S_1_L_4_out, I0 =>  inp_feat(11), I1 =>  inp_feat(508), I2 =>  inp_feat(466), I3 =>  inp_feat(41), I4 =>  inp_feat(426), I5 =>  inp_feat(459), I6 =>  inp_feat(477), I7 =>  inp_feat(143)); 
C_7_S_1_L_5_inst : LUT8 generic map(INIT => "1110010000100000000101000000010000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000011101100111101100001010001000100000000000000000000000000000000000100000001110101000001000101010100000000000000000000000000000000") port map( O =>C_7_S_1_L_5_out, I0 =>  inp_feat(366), I1 =>  inp_feat(427), I2 =>  inp_feat(290), I3 =>  inp_feat(486), I4 =>  inp_feat(311), I5 =>  inp_feat(328), I6 =>  inp_feat(411), I7 =>  inp_feat(170)); 
C_7_S_1_L_6_inst : LUT8 generic map(INIT => "0001001110110011000011010011011110010001000000011000000100100001000000000010000000000000000000000000000000000000000000000000000000000000000000010000000100000011000000010000000000000000000000100000000000000000000000000000001000000000000100000000000000000000") port map( O =>C_7_S_1_L_6_out, I0 =>  inp_feat(57), I1 =>  inp_feat(487), I2 =>  inp_feat(190), I3 =>  inp_feat(198), I4 =>  inp_feat(414), I5 =>  inp_feat(496), I6 =>  inp_feat(466), I7 =>  inp_feat(22)); 
C_7_S_1_L_7_inst : LUT8 generic map(INIT => "1010111010101110000010101010001000101000000011000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_1_L_7_out, I0 =>  inp_feat(280), I1 =>  inp_feat(151), I2 =>  inp_feat(98), I3 =>  inp_feat(65), I4 =>  inp_feat(444), I5 =>  inp_feat(183), I6 =>  inp_feat(325), I7 =>  inp_feat(212)); 
C_7_S_2_L_0_inst : LUT8 generic map(INIT => "0100100000000000001001001100010010001000000010000000000000000000000001000000000000000000010000000000000000000000000000000000000011000100110000000000010011000000000000000000100000000000000011000000010000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_2_L_0_out, I0 =>  inp_feat(190), I1 =>  inp_feat(15), I2 =>  inp_feat(382), I3 =>  inp_feat(350), I4 =>  inp_feat(446), I5 =>  inp_feat(459), I6 =>  inp_feat(143), I7 =>  inp_feat(503)); 
C_7_S_2_L_1_inst : LUT8 generic map(INIT => "1010000010001000000001000000000010000000000000000000000000000000111000001000000001001011000000101100000011000000000000000000000010000010000000000000000000000000000000000000000000000000000000001000000000000000010000100000000000000000000000000000000000000000") port map( O =>C_7_S_2_L_1_out, I0 =>  inp_feat(351), I1 =>  inp_feat(352), I2 =>  inp_feat(478), I3 =>  inp_feat(297), I4 =>  inp_feat(180), I5 =>  inp_feat(178), I6 =>  inp_feat(437), I7 =>  inp_feat(340)); 
C_7_S_2_L_2_inst : LUT8 generic map(INIT => "0101000111110100010000000001000011000000011001001100000000000000001000100001000000000000000000000000000000000000000000000000000001110001110100010101000101110010010000000000000000000000000001010000000000000000011100000101000000000000000000000000000000000000") port map( O =>C_7_S_2_L_2_out, I0 =>  inp_feat(503), I1 =>  inp_feat(290), I2 =>  inp_feat(374), I3 =>  inp_feat(258), I4 =>  inp_feat(212), I5 =>  inp_feat(496), I6 =>  inp_feat(466), I7 =>  inp_feat(440)); 
C_7_S_2_L_3_inst : LUT8 generic map(INIT => "1111100011010000110100000000000000000000110000000000000001000000000010000101000010001000010000000000000000010000000000000001000000000000000000000000000000000100000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_2_L_3_out, I0 =>  inp_feat(190), I1 =>  inp_feat(502), I2 =>  inp_feat(86), I3 =>  inp_feat(264), I4 =>  inp_feat(61), I5 =>  inp_feat(311), I6 =>  inp_feat(496), I7 =>  inp_feat(143)); 
C_7_S_2_L_4_inst : LUT8 generic map(INIT => "1000010010100000010000001010000010000000001010000000000000000000001100000000000000000000000000000000000000000000000000000000000010110001111100100000000000010100110111111111100110011101101100010000000000000000000000000000000010000100101100000000000001000000") port map( O =>C_7_S_2_L_4_out, I0 =>  inp_feat(496), I1 =>  inp_feat(350), I2 =>  inp_feat(224), I3 =>  inp_feat(100), I4 =>  inp_feat(112), I5 =>  inp_feat(166), I6 =>  inp_feat(466), I7 =>  inp_feat(422)); 
C_7_S_2_L_5_inst : LUT8 generic map(INIT => "1000001010000000111010000000000000000000000000001010100000000000000100101000000000000000000000000000000000000000000000000000000000000110000000000000010000000000000010001000000000010100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_2_L_5_out, I0 =>  inp_feat(373), I1 =>  inp_feat(80), I2 =>  inp_feat(120), I3 =>  inp_feat(327), I4 =>  inp_feat(171), I5 =>  inp_feat(459), I6 =>  inp_feat(306), I7 =>  inp_feat(374)); 
C_7_S_2_L_6_inst : LUT8 generic map(INIT => "1010000000000001000001100000000010000000000000001100000000000000101010001000000010001000000000001000000000000000010001000000000010000000000000000000000000000000000000000000000011000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_2_L_6_out, I0 =>  inp_feat(41), I1 =>  inp_feat(328), I2 =>  inp_feat(290), I3 =>  inp_feat(248), I4 =>  inp_feat(201), I5 =>  inp_feat(385), I6 =>  inp_feat(446), I7 =>  inp_feat(112)); 
C_7_S_2_L_7_inst : LUT8 generic map(INIT => "1010000010100000100000000000000000100000101000001000000000000000100000000000000011000000000000001000000000000000110000000000000000000000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_2_L_7_out, I0 =>  inp_feat(15), I1 =>  inp_feat(10), I2 =>  inp_feat(241), I3 =>  inp_feat(353), I4 =>  inp_feat(420), I5 =>  inp_feat(382), I6 =>  inp_feat(427), I7 =>  inp_feat(341)); 
C_7_S_3_L_0_inst : LUT8 generic map(INIT => "1100011101000001000100000000000011111111000100100000000000000000010001010010000000000000000100001111111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000") port map( O =>C_7_S_3_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(362), I2 =>  inp_feat(234), I3 =>  inp_feat(394), I4 =>  inp_feat(259), I5 =>  inp_feat(498), I6 =>  inp_feat(275), I7 =>  inp_feat(387)); 
C_7_S_3_L_1_inst : LUT8 generic map(INIT => "1010000010000000101010100000000000010000001000000000000000000000100000001100000000000100110000000000000000000000000000001100000000000000000000001000100100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_3_L_1_out, I0 =>  inp_feat(154), I1 =>  inp_feat(275), I2 =>  inp_feat(11), I3 =>  inp_feat(229), I4 =>  inp_feat(210), I5 =>  inp_feat(376), I6 =>  inp_feat(180), I7 =>  inp_feat(178)); 
C_7_S_3_L_2_inst : LUT8 generic map(INIT => "0000001000100000101000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000100100101000001010000000000000111000000000000000000000000000001110100000100000001000000000000000100000000000000000000000000000") port map( O =>C_7_S_3_L_2_out, I0 =>  inp_feat(459), I1 =>  inp_feat(378), I2 =>  inp_feat(15), I3 =>  inp_feat(353), I4 =>  inp_feat(70), I5 =>  inp_feat(471), I6 =>  inp_feat(61), I7 =>  inp_feat(347)); 
C_7_S_3_L_3_inst : LUT8 generic map(INIT => "0001110001010100010011001000111000000000000001110010000011100111000010000000000000000000000000000000000000000000000000100000010010000010001000000000000000000001000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_3_L_3_out, I0 =>  inp_feat(492), I1 =>  inp_feat(381), I2 =>  inp_feat(258), I3 =>  inp_feat(198), I4 =>  inp_feat(100), I5 =>  inp_feat(76), I6 =>  inp_feat(459), I7 =>  inp_feat(306)); 
C_7_S_3_L_4_inst : LUT8 generic map(INIT => "1000001000000000011111000000000000100000000000000100000000100010011110010000000011110000000000000000000000000000001001000000000010000000000000000000000000000000000000000000000000000000100000100010010000000000100000000000000000010000000000000000000000000000") port map( O =>C_7_S_3_L_4_out, I0 =>  inp_feat(98), I1 =>  inp_feat(100), I2 =>  inp_feat(478), I3 =>  inp_feat(116), I4 =>  inp_feat(331), I5 =>  inp_feat(480), I6 =>  inp_feat(382), I7 =>  inp_feat(212)); 
C_7_S_3_L_5_inst : LUT8 generic map(INIT => "0010000000000000000000001000000010111010010000100000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000000000000100010000000111011000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_7_S_3_L_5_out, I0 =>  inp_feat(451), I1 =>  inp_feat(13), I2 =>  inp_feat(467), I3 =>  inp_feat(321), I4 =>  inp_feat(365), I5 =>  inp_feat(362), I6 =>  inp_feat(266), I7 =>  inp_feat(382)); 
C_7_S_3_L_6_inst : LUT8 generic map(INIT => "1010001101110000101000000000000000000000000000000000000000000000110000101100000010001011000000000000000000000000000000000000000010000000001000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_3_L_6_out, I0 =>  inp_feat(154), I1 =>  inp_feat(336), I2 =>  inp_feat(204), I3 =>  inp_feat(478), I4 =>  inp_feat(11), I5 =>  inp_feat(266), I6 =>  inp_feat(446), I7 =>  inp_feat(112)); 
C_7_S_3_L_7_inst : LUT8 generic map(INIT => "1100100101010101010000000101001111000000011100000100010101010100110000000110001011000000011110010111001101101000010010001111111100000000000000000000000000000000100000000001000000000000001100000000010000000000000000000010100011110000000100000000010010011001") port map( O =>C_7_S_3_L_7_out, I0 =>  inp_feat(508), I1 =>  inp_feat(219), I2 =>  inp_feat(427), I3 =>  inp_feat(503), I4 =>  inp_feat(486), I5 =>  inp_feat(382), I6 =>  inp_feat(98), I7 =>  inp_feat(458)); 
C_7_S_4_L_0_inst : LUT8 generic map(INIT => "1000001010100110100000001000000000000000110000000010100010000000110000001100010000000000100000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000") port map( O =>C_7_S_4_L_0_out, I0 =>  inp_feat(502), I1 =>  inp_feat(307), I2 =>  inp_feat(109), I3 =>  inp_feat(65), I4 =>  inp_feat(401), I5 =>  inp_feat(416), I6 =>  inp_feat(79), I7 =>  inp_feat(277)); 
C_7_S_4_L_1_inst : LUT8 generic map(INIT => "0011000101000001000000000000000000100010000000000000000000000000110100011101000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010100000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_4_L_1_out, I0 =>  inp_feat(385), I1 =>  inp_feat(258), I2 =>  inp_feat(381), I3 =>  inp_feat(143), I4 =>  inp_feat(92), I5 =>  inp_feat(24), I6 =>  inp_feat(85), I7 =>  inp_feat(224)); 
C_7_S_4_L_2_inst : LUT8 generic map(INIT => "1101100010000000100010000000000000000000100000001000000011000000100000000000000000000000000000000000000000000000100000000000000000000000001010000000001000100000000000000000000010000000001000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_7_S_4_L_2_out, I0 =>  inp_feat(480), I1 =>  inp_feat(222), I2 =>  inp_feat(173), I3 =>  inp_feat(509), I4 =>  inp_feat(170), I5 =>  inp_feat(11), I6 =>  inp_feat(311), I7 =>  inp_feat(496)); 
C_7_S_4_L_3_inst : LUT8 generic map(INIT => "1100111000111100100000000001000001000101000101011000000000000000110010100100000000010000000000001100111000000110000000000000000001000000001000000000000000000000010100000000000000000000000000000000000001010000000000000000000000000001000000000000000000000000") port map( O =>C_7_S_4_L_3_out, I0 =>  inp_feat(57), I1 =>  inp_feat(496), I2 =>  inp_feat(100), I3 =>  inp_feat(61), I4 =>  inp_feat(484), I5 =>  inp_feat(85), I6 =>  inp_feat(446), I7 =>  inp_feat(112)); 
C_7_S_4_L_4_inst : LUT8 generic map(INIT => "1101010101110100101100000100000010100000000000000000000000000000001000000010001000000000010000000000000000000000000000000000000010000000000010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_4_L_4_out, I0 =>  inp_feat(355), I1 =>  inp_feat(331), I2 =>  inp_feat(448), I3 =>  inp_feat(232), I4 =>  inp_feat(180), I5 =>  inp_feat(178), I6 =>  inp_feat(297), I7 =>  inp_feat(340)); 
C_7_S_4_L_5_inst : LUT8 generic map(INIT => "1111010001110111101100100000000010010000000000000000000000000000000000001000100100000010000000000000000000000001000000000000000000000000010010100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_7_S_4_L_5_out, I0 =>  inp_feat(59), I1 =>  inp_feat(504), I2 =>  inp_feat(232), I3 =>  inp_feat(98), I4 =>  inp_feat(180), I5 =>  inp_feat(178), I6 =>  inp_feat(297), I7 =>  inp_feat(340)); 
C_7_S_4_L_6_inst : LUT8 generic map(INIT => "1000100010011000000000000000001000000011100001000000000000000000000000000000000000001000000000000000000000000000000000000000000011101110111001001110101101000010110110001010000000111100000000000100100001000000010001001000000000000000000000001110000000000000") port map( O =>C_7_S_4_L_6_out, I0 =>  inp_feat(434), I1 =>  inp_feat(381), I2 =>  inp_feat(22), I3 =>  inp_feat(224), I4 =>  inp_feat(76), I5 =>  inp_feat(458), I6 =>  inp_feat(288), I7 =>  inp_feat(198)); 
C_7_S_4_L_7_inst : LUT8 generic map(INIT => "1110000000000000000000001000000011110000100000001000000010000000000000000000000000000000000000000110000000000000000000000000000010010000101001000000000000000000100000000000000000000000000011001000000000000000000000000000000000000000000010000000000000000000") port map( O =>C_7_S_4_L_7_out, I0 =>  inp_feat(381), I1 =>  inp_feat(41), I2 =>  inp_feat(203), I3 =>  inp_feat(53), I4 =>  inp_feat(59), I5 =>  inp_feat(508), I6 =>  inp_feat(466), I7 =>  inp_feat(224)); 
C_8_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_0_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_1_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_2_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_3_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_8_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001000000010001000100010001000000000000000000000000000") port map( O =>C_8_S_4_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(5), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_0_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_0_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_1_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_1_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_2_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_2_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_3_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_3_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_9_S_4_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_9_S_4_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_10_S_0_L_0_inst : LUT8 generic map(INIT => "1111111010110000101110101011000010111000100000001011100010000000111110110010001110111011101100110000100000001000000010000000000011011000110100000011000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_10_S_0_L_0_out, I0 =>  inp_feat(51), I1 =>  inp_feat(212), I2 =>  inp_feat(280), I3 =>  inp_feat(398), I4 =>  inp_feat(411), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_10_S_0_L_1_inst : LUT8 generic map(INIT => "1010101010110011100000111011001100100111111100010000000110110001101010101110001000000000000000001000001011100010000000001100000010101010100000001000000010000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000") port map( O =>C_10_S_0_L_1_out, I0 =>  inp_feat(51), I1 =>  inp_feat(400), I2 =>  inp_feat(398), I3 =>  inp_feat(171), I4 =>  inp_feat(254), I5 =>  inp_feat(290), I6 =>  inp_feat(272), I7 =>  inp_feat(284)); 
C_10_S_0_L_2_inst : LUT8 generic map(INIT => "0010101001111111110110000000101010101010101010111010100000001000101000101010011100000010000000101000101100011111000000100000001110101010000011100000000000000000101010100000101100000000000000000000100000000110000000000000000000001011000011110000001000000010") port map( O =>C_10_S_0_L_2_out, I0 =>  inp_feat(398), I1 =>  inp_feat(405), I2 =>  inp_feat(323), I3 =>  inp_feat(224), I4 =>  inp_feat(477), I5 =>  inp_feat(289), I6 =>  inp_feat(311), I7 =>  inp_feat(100)); 
C_10_S_0_L_3_inst : LUT8 generic map(INIT => "1111110011110000111110000001000011111000000000000000000000000000111010000000000000000000000000000000000000000000000000000000000011011000000000000101100000000000110110000000000011110000000000000000000000000000000000000000000000001000000000000000000000000000") port map( O =>C_10_S_0_L_3_out, I0 =>  inp_feat(411), I1 =>  inp_feat(224), I2 =>  inp_feat(220), I3 =>  inp_feat(257), I4 =>  inp_feat(112), I5 =>  inp_feat(326), I6 =>  inp_feat(284), I7 =>  inp_feat(314)); 
C_10_S_0_L_4_inst : LUT8 generic map(INIT => "1111110011110000110111110001001011100111001000001110011100110010101000000010000000000000000000001010000000100000001000000010000011110001000100010000010101110001111111111111001101110111011001111000100010000000000000000000000011010101010001000101000100110101") port map( O =>C_10_S_0_L_4_out, I0 =>  inp_feat(487), I1 =>  inp_feat(496), I2 =>  inp_feat(292), I3 =>  inp_feat(398), I4 =>  inp_feat(102), I5 =>  inp_feat(212), I6 =>  inp_feat(51), I7 =>  inp_feat(446)); 
C_10_S_0_L_5_inst : LUT8 generic map(INIT => "1110000010101000010010000000000011100000101000001100100000000000111000001010000001001000000000001100100000000000100010000000000010000000000000001000100000000000100000000000000010001000000000000000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_10_S_0_L_5_out, I0 =>  inp_feat(257), I1 =>  inp_feat(424), I2 =>  inp_feat(284), I3 =>  inp_feat(220), I4 =>  inp_feat(311), I5 =>  inp_feat(411), I6 =>  inp_feat(466), I7 =>  inp_feat(22)); 
C_10_S_0_L_6_inst : LUT8 generic map(INIT => "1110100011001110001001001101100011100000101010001010100010100000000010101110000000000000111100000000000000000000001000000000000011101000111111101001000011110000000000001010101010100000101010000000000000100000000000000001000000000000000000000000000010000000") port map( O =>C_10_S_0_L_6_out, I0 =>  inp_feat(51), I1 =>  inp_feat(398), I2 =>  inp_feat(477), I3 =>  inp_feat(212), I4 =>  inp_feat(166), I5 =>  inp_feat(268), I6 =>  inp_feat(236), I7 =>  inp_feat(466)); 
C_10_S_0_L_7_inst : LUT8 generic map(INIT => "1010101101001111110011101100110011111111110000111010001000000010110000000101000000000010000000101110001001000010000000100000000011111111111000101000000000000000111110111100001000000000000000001111111001000010000000000000000001010010010000000000000000000000") port map( O =>C_10_S_0_L_7_out, I0 =>  inp_feat(57), I1 =>  inp_feat(374), I2 =>  inp_feat(458), I3 =>  inp_feat(398), I4 =>  inp_feat(184), I5 =>  inp_feat(306), I6 =>  inp_feat(317), I7 =>  inp_feat(378)); 
C_10_S_1_L_0_inst : LUT8 generic map(INIT => "1110110011101100100010001000100010101000101010000000100010001000111010101010100010000000100010001110000010001000000000000000100010100000101010001000000010001000101000001000100010001000100010001010101010101000000010001000100010101000100010000000100010001000") port map( O =>C_10_S_1_L_0_out, I0 =>  inp_feat(220), I1 =>  inp_feat(127), I2 =>  inp_feat(374), I3 =>  inp_feat(411), I4 =>  inp_feat(22), I5 =>  inp_feat(466), I6 =>  inp_feat(471), I7 =>  inp_feat(102)); 
C_10_S_1_L_1_inst : LUT8 generic map(INIT => "1111110011111000111100101111000011101000000000000010000000110000110011001110000000001000111100000000000000000000000000000000000010001000101010000000000010100000000000000000000000000000000000000000100000100000000000000010000000000000000000000000000000000000") port map( O =>C_10_S_1_L_1_out, I0 =>  inp_feat(459), I1 =>  inp_feat(200), I2 =>  inp_feat(430), I3 =>  inp_feat(38), I4 =>  inp_feat(272), I5 =>  inp_feat(284), I6 =>  inp_feat(370), I7 =>  inp_feat(352)); 
C_10_S_1_L_2_inst : LUT8 generic map(INIT => "1111011110111111101000111010101110101110101010001010000000000000100100000001011100000000000000000000001000001000000000000000000010110011101000111010000010000001001000000000000000000000000000000011000100110011000000000000000100000000000000000000000000000000") port map( O =>C_10_S_1_L_2_out, I0 =>  inp_feat(487), I1 =>  inp_feat(323), I2 =>  inp_feat(427), I3 =>  inp_feat(468), I4 =>  inp_feat(317), I5 =>  inp_feat(356), I6 =>  inp_feat(102), I7 =>  inp_feat(280)); 
C_10_S_1_L_3_inst : LUT8 generic map(INIT => "1010111010101110101010000000000010001100100000000000000000000000110111110001111100000000000000000000000000000000000000000000000011001100100011011110100000001000110011001000100010000000000000000101010101110011111000000000000000000000000000000000000000000000") port map( O =>C_10_S_1_L_3_out, I0 =>  inp_feat(137), I1 =>  inp_feat(458), I2 =>  inp_feat(496), I3 =>  inp_feat(102), I4 =>  inp_feat(199), I5 =>  inp_feat(352), I6 =>  inp_feat(326), I7 =>  inp_feat(143)); 
C_10_S_1_L_4_inst : LUT8 generic map(INIT => "0111110110100111111111100010011101111100011111010010011000100101111011101101111111101011111111110000101011111111000000100001011100001000100000001000100000100000101010000010000000001000001000001000100000000010101010000001001100000000001100000000000000100000") port map( O =>C_10_S_1_L_4_out, I0 =>  inp_feat(11), I1 =>  inp_feat(98), I2 =>  inp_feat(219), I3 =>  inp_feat(400), I4 =>  inp_feat(458), I5 =>  inp_feat(57), I6 =>  inp_feat(212), I7 =>  inp_feat(50)); 
C_10_S_1_L_5_inst : LUT8 generic map(INIT => "0111101111111111101111111001111111100010011011111000101100111111111100001111001011110011011100111010101000001110001100110011111110000110100001000001101110011011000010000000000000011010000001110000000000000000000100010101000100000000000000100001000000010111") port map( O =>C_10_S_1_L_5_out, I0 =>  inp_feat(468), I1 =>  inp_feat(289), I2 =>  inp_feat(137), I3 =>  inp_feat(458), I4 =>  inp_feat(400), I5 =>  inp_feat(76), I6 =>  inp_feat(276), I7 =>  inp_feat(398)); 
C_10_S_1_L_6_inst : LUT8 generic map(INIT => "1111110001010110011011000010101001001100000011111110110000000010101000000010001010100010001000100010001000000010000000000000001011100000111100001010111000100010000000000000001011001100000000101010000000100010101000100010001000000000000000000000000000000010") port map( O =>C_10_S_1_L_6_out, I0 =>  inp_feat(53), I1 =>  inp_feat(474), I2 =>  inp_feat(382), I3 =>  inp_feat(143), I4 =>  inp_feat(289), I5 =>  inp_feat(51), I6 =>  inp_feat(22), I7 =>  inp_feat(280)); 
C_10_S_1_L_7_inst : LUT8 generic map(INIT => "1111111111000000100000000000000011111100111100001000000000000000001100100000000000000000000000000011000000100000000000000000000000111010010000001000100000000000111010001100000010000000000000000000100000100000100000000000000010100000001000001000000000000000") port map( O =>C_10_S_1_L_7_out, I0 =>  inp_feat(102), I1 =>  inp_feat(143), I2 =>  inp_feat(51), I3 =>  inp_feat(501), I4 =>  inp_feat(284), I5 =>  inp_feat(452), I6 =>  inp_feat(199), I7 =>  inp_feat(88)); 
C_10_S_2_L_0_inst : LUT8 generic map(INIT => "1110100010000000111111111001111111110000100000001000000000000000111100000000000000000000000000000000000000000000000000000000000010110000000000001111011110001111000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_10_S_2_L_0_out, I0 =>  inp_feat(112), I1 =>  inp_feat(276), I2 =>  inp_feat(76), I3 =>  inp_feat(343), I4 =>  inp_feat(326), I5 =>  inp_feat(220), I6 =>  inp_feat(430), I7 =>  inp_feat(102)); 
C_10_S_2_L_1_inst : LUT8 generic map(INIT => "1110110011001000100011001100000011101100111011001101110100000100000000000100000010110100010000000001101000000000101010110000000000000000000000001000110000000000110111100100010010000111000000000000000000000000000011000000000000000010000000000010101000000000") port map( O =>C_10_S_2_L_1_out, I0 =>  inp_feat(468), I1 =>  inp_feat(236), I2 =>  inp_feat(60), I3 =>  inp_feat(50), I4 =>  inp_feat(121), I5 =>  inp_feat(400), I6 =>  inp_feat(430), I7 =>  inp_feat(102)); 
C_10_S_2_L_2_inst : LUT8 generic map(INIT => "1111001010100000101110101010001010111010100000000011001000100000111100000101000010110011001100111101000011000010001100110011000110111010101000001111101010000000000100000000000000001000000000000011011100010000111100010011000100010001000000001101001100010011") port map( O =>C_10_S_2_L_2_out, I0 =>  inp_feat(496), I1 =>  inp_feat(212), I2 =>  inp_feat(51), I3 =>  inp_feat(50), I4 =>  inp_feat(405), I5 =>  inp_feat(398), I6 =>  inp_feat(400), I7 =>  inp_feat(468)); 
C_10_S_2_L_3_inst : LUT8 generic map(INIT => "1110000000010000111111101100100000000000000000001000101000001000111110000111100010001010001010100010100000000000000010100000101011001100110000001100111011001010000011000000000000001110000000101000100000000000100010001010100000001000000000000000001000001010") port map( O =>C_10_S_2_L_3_out, I0 =>  inp_feat(494), I1 =>  inp_feat(50), I2 =>  inp_feat(377), I3 =>  inp_feat(398), I4 =>  inp_feat(212), I5 =>  inp_feat(76), I6 =>  inp_feat(292), I7 =>  inp_feat(85)); 
C_10_S_2_L_4_inst : LUT8 generic map(INIT => "0101110111011100111001011101000011001100110110001101100001010000100001000000000000000000010000001100110000000000000010000000000011001101100010000100010000000000110011001000010010000100000001001100000011001000100000000000010011001100110001001100110000000100") port map( O =>C_10_S_2_L_4_out, I0 =>  inp_feat(400), I1 =>  inp_feat(236), I2 =>  inp_feat(468), I3 =>  inp_feat(50), I4 =>  inp_feat(398), I5 =>  inp_feat(458), I6 =>  inp_feat(124), I7 =>  inp_feat(405)); 
C_10_S_2_L_5_inst : LUT8 generic map(INIT => "1110110001110101110011001000110011010001011101011111000011010100110011000000010100000000000000010000000100010101010000000001011100110001011100000100010000010001001101000011010111010100001100001001110101010101000001010000000001111100000101000111110000010001") port map( O =>C_10_S_2_L_5_out, I0 =>  inp_feat(323), I1 =>  inp_feat(98), I2 =>  inp_feat(288), I3 =>  inp_feat(487), I4 =>  inp_feat(166), I5 =>  inp_feat(382), I6 =>  inp_feat(143), I7 =>  inp_feat(224)); 
C_10_S_2_L_6_inst : LUT8 generic map(INIT => "1111100000011010111110011010111111011001100010101111111111111111111110001011101111111110101111110000000000010011010001010101011101001000000010000000100000001010000000000000000011011001100110011100100000111000101110010000101100000100000100000000000000010011") port map( O =>C_10_S_2_L_6_out, I0 =>  inp_feat(292), I1 =>  inp_feat(426), I2 =>  inp_feat(112), I3 =>  inp_feat(76), I4 =>  inp_feat(289), I5 =>  inp_feat(276), I6 =>  inp_feat(101), I7 =>  inp_feat(398)); 
C_10_S_2_L_7_inst : LUT8 generic map(INIT => "1011000011110010101000000010000010101010000000001000000000000000111100001111000000000000000000001000000000000000000000000000000010101000111010101100000011101010101010000000000000000000000000000000000011000000000000000000000010100000000000000000000000000000") port map( O =>C_10_S_2_L_7_out, I0 =>  inp_feat(199), I1 =>  inp_feat(366), I2 =>  inp_feat(102), I3 =>  inp_feat(143), I4 =>  inp_feat(51), I5 =>  inp_feat(388), I6 =>  inp_feat(262), I7 =>  inp_feat(400)); 
C_10_S_3_L_0_inst : LUT8 generic map(INIT => "0010111010101010101000110010100011111101011011110010000100000000111000001100000010100000000000000000000000000000000000000000000011101111110111001010011100000011111111110100111100100011000000011110000011000000101000000000000010000000000000001010000000000000") port map( O =>C_10_S_3_L_0_out, I0 =>  inp_feat(102), I1 =>  inp_feat(50), I2 =>  inp_feat(459), I3 =>  inp_feat(398), I4 =>  inp_feat(14), I5 =>  inp_feat(112), I6 =>  inp_feat(346), I7 =>  inp_feat(411)); 
C_10_S_3_L_1_inst : LUT8 generic map(INIT => "0010111011101100101001001000000011001100110011001000000010000000100010000000110000000000000000001100100000001100110010000000000011101010111011101000000000000000100011001000100010001000000000000000100010001000000000000000000010001000100010001000100000000000") port map( O =>C_10_S_3_L_1_out, I0 =>  inp_feat(398), I1 =>  inp_feat(111), I2 =>  inp_feat(190), I3 =>  inp_feat(311), I4 =>  inp_feat(177), I5 =>  inp_feat(170), I6 =>  inp_feat(258), I7 =>  inp_feat(378)); 
C_10_S_3_L_2_inst : LUT8 generic map(INIT => "1101110011000101000001001000010111100100100000000000000000100000111111001100010010100100110001000000000000000000000000000000000011101110100001001010110011000101001000001000000000000000100000001110111011000100101000001100010000000000000000000000000000000000") port map( O =>C_10_S_3_L_2_out, I0 =>  inp_feat(426), I1 =>  inp_feat(398), I2 =>  inp_feat(76), I3 =>  inp_feat(55), I4 =>  inp_feat(317), I5 =>  inp_feat(360), I6 =>  inp_feat(190), I7 =>  inp_feat(378)); 
C_10_S_3_L_3_inst : LUT8 generic map(INIT => "1110111001111101101000001110010111000000110000000000000000000000011101101110011100000001101001011100000011000000000000000000000010101111010001000010000001100100000000000000000000000000000000001100010001000100000000000000000011000000000000000000000000000000") port map( O =>C_10_S_3_L_3_out, I0 =>  inp_feat(68), I1 =>  inp_feat(166), I2 =>  inp_feat(22), I3 =>  inp_feat(340), I4 =>  inp_feat(51), I5 =>  inp_feat(263), I6 =>  inp_feat(224), I7 =>  inp_feat(477)); 
C_10_S_3_L_4_inst : LUT8 generic map(INIT => "0011110000110000010010000111000011011000011100001111100010010000111111001111000011001000101000001101100011110000110110001111000011111000111100001010000001110000111110001011000011111000111100000000000011110000000000001011000000000000101100001000000011110000") port map( O =>C_10_S_3_L_4_out, I0 =>  inp_feat(276), I1 =>  inp_feat(112), I2 =>  inp_feat(287), I3 =>  inp_feat(288), I4 =>  inp_feat(496), I5 =>  inp_feat(468), I6 =>  inp_feat(378), I7 =>  inp_feat(466)); 
C_10_S_3_L_5_inst : LUT8 generic map(INIT => "0100111111111101000111101000000010101011101010101000101110000000110000011111000001000001000000000000000100000000000000000000000011111111110111011101110100000000110111111001111100001001000001010000010100000000000000010000000000000001000000010000000000000000") port map( O =>C_10_S_3_L_5_out, I0 =>  inp_feat(98), I1 =>  inp_feat(102), I2 =>  inp_feat(233), I3 =>  inp_feat(385), I4 =>  inp_feat(398), I5 =>  inp_feat(219), I6 =>  inp_feat(184), I7 =>  inp_feat(411)); 
C_10_S_3_L_6_inst : LUT8 generic map(INIT => "1111000011101000111000010111000011010000000000000000000000000000111111011111110101010000111111011000000000000000000100000001000000000000111100000000000010001000101010001000000010000000000000001101010111011110111100001101010100000000000000001101101101110001") port map( O =>C_10_S_3_L_6_out, I0 =>  inp_feat(289), I1 =>  inp_feat(276), I2 =>  inp_feat(398), I3 =>  inp_feat(112), I4 =>  inp_feat(76), I5 =>  inp_feat(55), I6 =>  inp_feat(400), I7 =>  inp_feat(50)); 
C_10_S_3_L_7_inst : LUT8 generic map(INIT => "1110110010000000101010000000000011001100110000001100000000000000101010101000000011101010000000000000000000000000000000000000000011001000010000001100100000000000110000001100000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_10_S_3_L_7_out, I0 =>  inp_feat(88), I1 =>  inp_feat(67), I2 =>  inp_feat(272), I3 =>  inp_feat(284), I4 =>  inp_feat(499), I5 =>  inp_feat(311), I6 =>  inp_feat(258), I7 =>  inp_feat(505)); 
C_10_S_4_L_0_inst : LUT8 generic map(INIT => "1110101011101000111110000000000011101100110000001111101111010101000010001000000011001100110101000100010011000000000000001100010111001111110100001000000011010001110001001101000011001101110111011100010111010101010001011101010101000001010001000000010111010101") port map( O =>C_10_S_4_L_0_out, I0 =>  inp_feat(370), I1 =>  inp_feat(422), I2 =>  inp_feat(224), I3 =>  inp_feat(289), I4 =>  inp_feat(405), I5 =>  inp_feat(268), I6 =>  inp_feat(374), I7 =>  inp_feat(212)); 
C_10_S_4_L_1_inst : LUT8 generic map(INIT => "0111100011111010111010101110000011111100110000000011110000000000001110100100000001101111000000000100011000000000001010100000000000001000000000001100110000000000000000000000000000001000000000000000111100000000000011110000000000001110000000000000010000000000") port map( O =>C_10_S_4_L_1_out, I0 =>  inp_feat(458), I1 =>  inp_feat(287), I2 =>  inp_feat(320), I3 =>  inp_feat(81), I4 =>  inp_feat(452), I5 =>  inp_feat(93), I6 =>  inp_feat(477), I7 =>  inp_feat(50)); 
C_10_S_4_L_2_inst : LUT8 generic map(INIT => "0000110010101100100000001010000010010101100011001000000010100000100110001000000010000000101000001110110000000000101000000000000011111101100010001000000011100000111011001000100010100000000000001111110000000000101000001000000011111101000000001010000000000000") port map( O =>C_10_S_4_L_2_out, I0 =>  inp_feat(76), I1 =>  inp_feat(398), I2 =>  inp_feat(343), I3 =>  inp_feat(89), I4 =>  inp_feat(494), I5 =>  inp_feat(468), I6 =>  inp_feat(496), I7 =>  inp_feat(411)); 
C_10_S_4_L_3_inst : LUT8 generic map(INIT => "1111110110101100110001001000000011111111001010000100010100000100111101010100000011000100000000000100011000000000000001010000000011110101101011000000010010000100000100100000000000000000000000000100010000000100000001000000010000000000000000000000000000000000") port map( O =>C_10_S_4_L_3_out, I0 =>  inp_feat(496), I1 =>  inp_feat(102), I2 =>  inp_feat(170), I3 =>  inp_feat(177), I4 =>  inp_feat(328), I5 =>  inp_feat(100), I6 =>  inp_feat(398), I7 =>  inp_feat(477)); 
C_10_S_4_L_4_inst : LUT8 generic map(INIT => "1111000000000100111100111110000100001000000000001111100000000000111011001111010011111110111111111000000000000000001100000000000011101110000000000100111001000111101000000000000000100000000000001110101010000010111111101111111111100000000000001010000000000000") port map( O =>C_10_S_4_L_4_out, I0 =>  inp_feat(290), I1 =>  inp_feat(493), I2 =>  inp_feat(326), I3 =>  inp_feat(137), I4 =>  inp_feat(191), I5 =>  inp_feat(134), I6 =>  inp_feat(190), I7 =>  inp_feat(378)); 
C_10_S_4_L_5_inst : LUT8 generic map(INIT => "1111001101110000110000001110000011111000000000000000000000000000111000000000000000000000000000000111000000000000000000000000000010101011001000000000000000000000111110100000000000000000000000001000000000000000000000000000000011111010000000000000000000000000") port map( O =>C_10_S_4_L_5_out, I0 =>  inp_feat(458), I1 =>  inp_feat(378), I2 =>  inp_feat(199), I3 =>  inp_feat(220), I4 =>  inp_feat(383), I5 =>  inp_feat(232), I6 =>  inp_feat(102), I7 =>  inp_feat(143)); 
C_10_S_4_L_6_inst : LUT8 generic map(INIT => "1010101011111011101100101010101000101000111100000010000000100000001010101010111110110010111011111010000000100000000100001010000010101010001000000011000010110000000000000000000001110000101000001010101000100000111100001011000000000000000000000011000010100000") port map( O =>C_10_S_4_L_6_out, I0 =>  inp_feat(51), I1 =>  inp_feat(212), I2 =>  inp_feat(437), I3 =>  inp_feat(468), I4 =>  inp_feat(374), I5 =>  inp_feat(398), I6 =>  inp_feat(458), I7 =>  inp_feat(22)); 
C_10_S_4_L_7_inst : LUT8 generic map(INIT => "0111101011001000111111110000000011111010110000001111001100000000111011001100110011001110110001001111001111001100011101111100110011000000110000001111010110000000010000000000000011110001100000001100010011000100000001001000000000100100110010000000010010000100") port map( O =>C_10_S_4_L_7_out, I0 =>  inp_feat(493), I1 =>  inp_feat(336), I2 =>  inp_feat(102), I3 =>  inp_feat(311), I4 =>  inp_feat(98), I5 =>  inp_feat(143), I6 =>  inp_feat(233), I7 =>  inp_feat(398)); 
C_11_S_0_L_0_inst : LUT8 generic map(INIT => "1110101111111010101010101110000010000000101000001010000010100000110000100000001010000000000000000000000000100000101000001010000011100010111000101010100011100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_0_out, I0 =>  inp_feat(507), I1 =>  inp_feat(291), I2 =>  inp_feat(238), I3 =>  inp_feat(472), I4 =>  inp_feat(378), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_11_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111101111101000110011111111101100000000000010000000100000110100011110101100000000000000100000000000000000000000000000000011101000110000000000000000000000100010000000000000000000000000001100000011000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(40), I2 =>  inp_feat(434), I3 =>  inp_feat(346), I4 =>  inp_feat(199), I5 =>  inp_feat(326), I6 =>  inp_feat(352), I7 =>  inp_feat(147)); 
C_11_S_0_L_2_inst : LUT8 generic map(INIT => "1111110010010010111000001010000001000000001100001110000011100000111011001000110011000000000000001100100000001000110000000000000011111100100000001010000010101000100000001000100010100000101000000000110000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_2_out, I0 =>  inp_feat(74), I1 =>  inp_feat(397), I2 =>  inp_feat(51), I3 =>  inp_feat(370), I4 =>  inp_feat(502), I5 =>  inp_feat(408), I6 =>  inp_feat(420), I7 =>  inp_feat(327)); 
C_11_S_0_L_3_inst : LUT8 generic map(INIT => "1000101011101010101010101011101111101110100010001010101110000100111010101110000010100010101000101000000000000000000000000000000011110100111111101000101011101011111101001100110000001100110010001100000001000000100000000010000010000000000000000000000000000000") port map( O =>C_11_S_0_L_3_out, I0 =>  inp_feat(370), I1 =>  inp_feat(291), I2 =>  inp_feat(457), I3 =>  inp_feat(492), I4 =>  inp_feat(399), I5 =>  inp_feat(302), I6 =>  inp_feat(385), I7 =>  inp_feat(6)); 
C_11_S_0_L_4_inst : LUT8 generic map(INIT => "1111110010001000111111110001000011110000111000001011000010110000010100000000000000110011001100000000000010110000001100001011000011000100000000001101110000000000110100001100000000000000000000000101000001000000011101010000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_4_out, I0 =>  inp_feat(195), I1 =>  inp_feat(496), I2 =>  inp_feat(352), I3 =>  inp_feat(350), I4 =>  inp_feat(382), I5 =>  inp_feat(327), I6 =>  inp_feat(398), I7 =>  inp_feat(428)); 
C_11_S_0_L_5_inst : LUT8 generic map(INIT => "1111110110111101111111001011110111000000101011101111010010100000100100000000000000000000001000000000000000000000000000000010000010101000100000001100100010000000100000001000000011010000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_5_out, I0 =>  inp_feat(64), I1 =>  inp_feat(474), I2 =>  inp_feat(131), I3 =>  inp_feat(327), I4 =>  inp_feat(6), I5 =>  inp_feat(41), I6 =>  inp_feat(67), I7 =>  inp_feat(19)); 
C_11_S_0_L_6_inst : LUT8 generic map(INIT => "1111111100101000111010001100100011111000101010001110100011001000100011100000000010001000000000000000000000000000000000000000000011111110100000001100100011000000111000001000000011000000110000000001111100000000100010000000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_6_out, I0 =>  inp_feat(324), I1 =>  inp_feat(134), I2 =>  inp_feat(382), I3 =>  inp_feat(326), I4 =>  inp_feat(327), I5 =>  inp_feat(366), I6 =>  inp_feat(19), I7 =>  inp_feat(304)); 
C_11_S_0_L_7_inst : LUT8 generic map(INIT => "1111110111110101111111111111111111001100101001001110110011101100111011000000000010000000100000000000000000000000100000000000000001010100010000000000010001000100010011000000010001000100010001001100110000000000100000000000000000000000000000000000000000000000") port map( O =>C_11_S_0_L_7_out, I0 =>  inp_feat(399), I1 =>  inp_feat(350), I2 =>  inp_feat(283), I3 =>  inp_feat(244), I4 =>  inp_feat(61), I5 =>  inp_feat(398), I6 =>  inp_feat(155), I7 =>  inp_feat(352)); 
C_11_S_1_L_0_inst : LUT8 generic map(INIT => "1110101111111010101010101110000010000000101000001010000010100000110000100000001010000000000000000000000000100000101000001010000011100010111000101010100011100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_1_L_0_out, I0 =>  inp_feat(507), I1 =>  inp_feat(291), I2 =>  inp_feat(238), I3 =>  inp_feat(472), I4 =>  inp_feat(378), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_11_S_1_L_1_inst : LUT8 generic map(INIT => "1111111111101111101000110011111111101100000000000010000000100000110100011110101100000000000000100000000000000000000000000000000011101000110000000000000000000000100010000000000000000000000000001100000011000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_1_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(40), I2 =>  inp_feat(434), I3 =>  inp_feat(346), I4 =>  inp_feat(199), I5 =>  inp_feat(326), I6 =>  inp_feat(352), I7 =>  inp_feat(147)); 
C_11_S_1_L_2_inst : LUT8 generic map(INIT => "1110100010100000111001000000000000100010100000000010000000000000111011101010100000001100000010001000111010001010000010000000100010101000101010001110000000000000101010000000000010100000000000001000000010100000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_1_L_2_out, I0 =>  inp_feat(199), I1 =>  inp_feat(362), I2 =>  inp_feat(434), I3 =>  inp_feat(416), I4 =>  inp_feat(317), I5 =>  inp_feat(408), I6 =>  inp_feat(420), I7 =>  inp_feat(327)); 
C_11_S_1_L_3_inst : LUT8 generic map(INIT => "1110100000000100110011000000100000000000000001000101100000001100111010000000010011101000110011001110100000000000111010000100110011100000000000001100000000000000110000000000000011000000000000001010000000000000000000000000000010000000000000000000000000000000") port map( O =>C_11_S_1_L_3_out, I0 =>  inp_feat(436), I1 =>  inp_feat(199), I2 =>  inp_feat(339), I3 =>  inp_feat(255), I4 =>  inp_feat(105), I5 =>  inp_feat(408), I6 =>  inp_feat(6), I7 =>  inp_feat(366)); 
C_11_S_1_L_4_inst : LUT8 generic map(INIT => "1111101011101000111110101010101011110001000000001111000000000000111110111000101001010000000000001111000101000000000000000000000000100000000000000101000010000000000000000000000000000000000000001100100010001000010000000000000000000000000000000000000000000000") port map( O =>C_11_S_1_L_4_out, I0 =>  inp_feat(145), I1 =>  inp_feat(88), I2 =>  inp_feat(398), I3 =>  inp_feat(100), I4 =>  inp_feat(327), I5 =>  inp_feat(240), I6 =>  inp_feat(121), I7 =>  inp_feat(489)); 
C_11_S_1_L_5_inst : LUT8 generic map(INIT => "1110111010101100111010001010100010101010101000001010101010101000110010000010100000000000001000000010000000100000000000001010000011001000000011001000000010000000001100000000000000000000100010000000100000001000000000000000000000000000000000000000000010000000") port map( O =>C_11_S_1_L_5_out, I0 =>  inp_feat(318), I1 =>  inp_feat(131), I2 =>  inp_feat(427), I3 =>  inp_feat(100), I4 =>  inp_feat(237), I5 =>  inp_feat(197), I6 =>  inp_feat(507), I7 =>  inp_feat(317)); 
C_11_S_1_L_6_inst : LUT8 generic map(INIT => "1110110010001000110011001100110010101010100000001000111110001111110000000000000011001000100000001000101000000000100011111000111110001000000010001000101010000000000000000000000010000000100000001000100000000000100010000000000010001000000010001000100010001000") port map( O =>C_11_S_1_L_6_out, I0 =>  inp_feat(342), I1 =>  inp_feat(489), I2 =>  inp_feat(297), I3 =>  inp_feat(428), I4 =>  inp_feat(224), I5 =>  inp_feat(434), I6 =>  inp_feat(244), I7 =>  inp_feat(370)); 
C_11_S_1_L_7_inst : LUT8 generic map(INIT => "1100100010001100110010001010101011001000100010001100100000000000010010001000000011001000100000001000100000000000110010000000000011111100110011001000100010001000110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_1_L_7_out, I0 =>  inp_feat(134), I1 =>  inp_feat(67), I2 =>  inp_feat(338), I3 =>  inp_feat(6), I4 =>  inp_feat(327), I5 =>  inp_feat(433), I6 =>  inp_feat(350), I7 =>  inp_feat(220)); 
C_11_S_2_L_0_inst : LUT8 generic map(INIT => "1110101111111010101010101110000010000000101000001010000010100000110000100000001010000000000000000000000000100000101000001010000011100010111000101010100011100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_2_L_0_out, I0 =>  inp_feat(507), I1 =>  inp_feat(291), I2 =>  inp_feat(238), I3 =>  inp_feat(472), I4 =>  inp_feat(378), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_11_S_2_L_1_inst : LUT8 generic map(INIT => "1111111111101111101000110011111111101100000000000010000000100000110100011110101100000000000000100000000000000000000000000000000011101000110000000000000000000000100010000000000000000000000000001100000011000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_2_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(40), I2 =>  inp_feat(434), I3 =>  inp_feat(346), I4 =>  inp_feat(199), I5 =>  inp_feat(326), I6 =>  inp_feat(352), I7 =>  inp_feat(147)); 
C_11_S_2_L_2_inst : LUT8 generic map(INIT => "1111101110101010111110000000000001110000010000000011000000000000111110101110101011110000110000001100000011000000111000001010000010111000101010001000000000000000101100000000000010000000000000001000000010100000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_2_L_2_out, I0 =>  inp_feat(285), I1 =>  inp_feat(362), I2 =>  inp_feat(433), I3 =>  inp_feat(416), I4 =>  inp_feat(391), I5 =>  inp_feat(408), I6 =>  inp_feat(420), I7 =>  inp_feat(327)); 
C_11_S_2_L_3_inst : LUT8 generic map(INIT => "1111101011111000110000000000000011100000110000000000000000000000010000001100000000000000000000001100000011001100000000000000000011101010110010001100000000000000101000001100000000000000000000001100000001000000000000000000000011000000110011000000000000000000") port map( O =>C_11_S_2_L_3_out, I0 =>  inp_feat(244), I1 =>  inp_feat(210), I2 =>  inp_feat(449), I3 =>  inp_feat(0), I4 =>  inp_feat(313), I5 =>  inp_feat(309), I6 =>  inp_feat(398), I7 =>  inp_feat(6)); 
C_11_S_2_L_4_inst : LUT8 generic map(INIT => "1111110111011101111110000000000010001000111111011000000000001000111100001100110011111100000000000000000000000000000000000000000011101000000101001000000000000000101010101100110100000000000000001000000011001100110011000000000000000000110011000000000000000000") port map( O =>C_11_S_2_L_4_out, I0 =>  inp_feat(318), I1 =>  inp_feat(419), I2 =>  inp_feat(290), I3 =>  inp_feat(310), I4 =>  inp_feat(326), I5 =>  inp_feat(87), I6 =>  inp_feat(244), I7 =>  inp_feat(100)); 
C_11_S_2_L_5_inst : LUT8 generic map(INIT => "1000110011101100111101001110110010110000101000001111000010100000101001001010010011000000110001001010000010100000101000000010000011100100100000000100010000000000111000001000000011110000000000001010000000000000000000000000000010100000000000000000000000000000") port map( O =>C_11_S_2_L_5_out, I0 =>  inp_feat(100), I1 =>  inp_feat(326), I2 =>  inp_feat(62), I3 =>  inp_feat(56), I4 =>  inp_feat(405), I5 =>  inp_feat(244), I6 =>  inp_feat(216), I7 =>  inp_feat(170)); 
C_11_S_2_L_6_inst : LUT8 generic map(INIT => "1011100010101010101110101010101011110011111111110111000000010000111100001011101010100010101100100111000000110000000000000010000000010000000000001001001010001010000000000000000000000000000000001111000010100010101000101010001010000000101000000000000000000000") port map( O =>C_11_S_2_L_6_out, I0 =>  inp_feat(110), I1 =>  inp_feat(323), I2 =>  inp_feat(398), I3 =>  inp_feat(6), I4 =>  inp_feat(436), I5 =>  inp_feat(370), I6 =>  inp_feat(81), I7 =>  inp_feat(416)); 
C_11_S_2_L_7_inst : LUT8 generic map(INIT => "1111111111111100011110001111110011111111111100001111000011110000111111001111010001000000111000001111111111110000000000001110000011001100110011000000000011000100110000000000000000000000000000000100110000000000000000000000000011000000100000000000000000000000") port map( O =>C_11_S_2_L_7_out, I0 =>  inp_feat(6), I1 =>  inp_feat(268), I2 =>  inp_feat(358), I3 =>  inp_feat(301), I4 =>  inp_feat(370), I5 =>  inp_feat(327), I6 =>  inp_feat(149), I7 =>  inp_feat(416)); 
C_11_S_3_L_0_inst : LUT8 generic map(INIT => "1110101111111010101010101110000010000000101000001010000010100000110000100000001010000000000000000000000000100000101000001010000011100010111000101010100011100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_3_L_0_out, I0 =>  inp_feat(507), I1 =>  inp_feat(291), I2 =>  inp_feat(238), I3 =>  inp_feat(472), I4 =>  inp_feat(378), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_11_S_3_L_1_inst : LUT8 generic map(INIT => "1111110111111111101000110011011111111100000000000010000000100000110100011111111100000000000000100000000000000000000000000000000011010100110000000000000000000000000001000000000000000000000000001100000011000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_3_L_1_out, I0 =>  inp_feat(427), I1 =>  inp_feat(40), I2 =>  inp_feat(434), I3 =>  inp_feat(346), I4 =>  inp_feat(199), I5 =>  inp_feat(326), I6 =>  inp_feat(352), I7 =>  inp_feat(147)); 
C_11_S_3_L_2_inst : LUT8 generic map(INIT => "1100110011001100110010001100000010101010000010000000000000001000100010001100100000000000100000001000100011001100000000000000100011001000100010000000100000000000100000000000100000000000000000001100000011001100000000000000000000000000100011000000000000000000") port map( O =>C_11_S_3_L_2_out, I0 =>  inp_feat(147), I1 =>  inp_feat(313), I2 =>  inp_feat(15), I3 =>  inp_feat(400), I4 =>  inp_feat(443), I5 =>  inp_feat(328), I6 =>  inp_feat(398), I7 =>  inp_feat(290)); 
C_11_S_3_L_3_inst : LUT8 generic map(INIT => "1110110011000000111000001100000011111000110000001110100010100000011100000100000011110000110000001111000000000000111110001010100011101000111000001100101000000000000000000000000010001000000000000000000011000000101010100000000000000000000000001010100010000000") port map( O =>C_11_S_3_L_3_out, I0 =>  inp_feat(385), I1 =>  inp_feat(265), I2 =>  inp_feat(199), I3 =>  inp_feat(51), I4 =>  inp_feat(400), I5 =>  inp_feat(413), I6 =>  inp_feat(422), I7 =>  inp_feat(505)); 
C_11_S_3_L_4_inst : LUT8 generic map(INIT => "1100111010001000110011001000100010100000000000001100110000000000110111001100000011001100100000001100000001000000110000000000000011110000110100000100000000000000111100000001000000000000000000001100000001010000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_3_L_4_out, I0 =>  inp_feat(323), I1 =>  inp_feat(489), I2 =>  inp_feat(220), I3 =>  inp_feat(398), I4 =>  inp_feat(331), I5 =>  inp_feat(507), I6 =>  inp_feat(293), I7 =>  inp_feat(434)); 
C_11_S_3_L_5_inst : LUT8 generic map(INIT => "1101000011111100111111001111110011111000101100001111001000100000110010001101000011000000110110001100110010000000100000001000000011110000000000001101000000000000110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_3_L_5_out, I0 =>  inp_feat(301), I1 =>  inp_feat(370), I2 =>  inp_feat(489), I3 =>  inp_feat(290), I4 =>  inp_feat(6), I5 =>  inp_feat(327), I6 =>  inp_feat(210), I7 =>  inp_feat(199)); 
C_11_S_3_L_6_inst : LUT8 generic map(INIT => "1111110011111100110010001000100010001000000000001001000000000000101010001110110000000000000000001000110010001000000000000000000011100000100000001101000000000000110100000000000011010000000000001100100011101000111100000000000011011000100010000111000000000000") port map( O =>C_11_S_3_L_6_out, I0 =>  inp_feat(370), I1 =>  inp_feat(350), I2 =>  inp_feat(84), I3 =>  inp_feat(81), I4 =>  inp_feat(164), I5 =>  inp_feat(398), I6 =>  inp_feat(434), I7 =>  inp_feat(244)); 
C_11_S_3_L_7_inst : LUT8 generic map(INIT => "1111101010111010111110000011000010101000000000001111100000001000101010001000100010110000001000000000000000100000000000001000000011000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_3_L_7_out, I0 =>  inp_feat(370), I1 =>  inp_feat(264), I2 =>  inp_feat(501), I3 =>  inp_feat(398), I4 =>  inp_feat(10), I5 =>  inp_feat(199), I6 =>  inp_feat(436), I7 =>  inp_feat(210)); 
C_11_S_4_L_0_inst : LUT8 generic map(INIT => "1110101111111010101010101110000010000000101000001010000010100000110000100000001010000000000000000000000000100000101000001010000011100010111000101010100011100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_4_L_0_out, I0 =>  inp_feat(507), I1 =>  inp_feat(291), I2 =>  inp_feat(238), I3 =>  inp_feat(472), I4 =>  inp_feat(378), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_11_S_4_L_1_inst : LUT8 generic map(INIT => "1110111011101111101000100010101010101100000000000010000000100000101000101010101100000000000000100000000000000000000000000000000010101000100000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_11_S_4_L_1_out, I0 =>  inp_feat(489), I1 =>  inp_feat(40), I2 =>  inp_feat(434), I3 =>  inp_feat(346), I4 =>  inp_feat(199), I5 =>  inp_feat(326), I6 =>  inp_feat(352), I7 =>  inp_feat(147)); 
C_11_S_4_L_2_inst : LUT8 generic map(INIT => "1111100011010000000010000000000011010000100000000000000000000000110110001100000010001000000000001101000000000000000000000000000011001100110000001100100010001000010000000000000011000000000000001101111011000000110010001000100011000000000000000000000000000000") port map( O =>C_11_S_4_L_2_out, I0 =>  inp_feat(143), I1 =>  inp_feat(199), I2 =>  inp_feat(449), I3 =>  inp_feat(352), I4 =>  inp_feat(62), I5 =>  inp_feat(350), I6 =>  inp_feat(6), I7 =>  inp_feat(100)); 
C_11_S_4_L_3_inst : LUT8 generic map(INIT => "1111111110101110000000001010000010101111000011110000000000000000001000010010000000000000000000000011011100011111000000000000000011110011111010101010000010100000001000110010111100000000000000001110000011100000000000000000000000100101001111110000000000000000") port map( O =>C_11_S_4_L_3_out, I0 =>  inp_feat(290), I1 =>  inp_feat(195), I2 =>  inp_feat(407), I3 =>  inp_feat(143), I4 =>  inp_feat(313), I5 =>  inp_feat(309), I6 =>  inp_feat(398), I7 =>  inp_feat(244)); 
C_11_S_4_L_4_inst : LUT8 generic map(INIT => "0111000111000000110110000000000011000000100000001101000000000000110010001100000010001000000000001100000010000000010000000000000011111011100010001000100000000000110100010000000010000000000000001000100000000000100010000000000000000000000000000000000000000000") port map( O =>C_11_S_4_L_4_out, I0 =>  inp_feat(273), I1 =>  inp_feat(199), I2 =>  inp_feat(350), I3 =>  inp_feat(424), I4 =>  inp_feat(382), I5 =>  inp_feat(375), I6 =>  inp_feat(487), I7 =>  inp_feat(327)); 
C_11_S_4_L_5_inst : LUT8 generic map(INIT => "1110111011101110111001001110111011001000010000001000000000000000111011111000100001000000000010001000100000000000000000000000000011011101100011001101011100000101100010000000000000000000000000000100011110001001000001110000010010001000000000000000000000000000") port map( O =>C_11_S_4_L_5_out, I0 =>  inp_feat(399), I1 =>  inp_feat(51), I2 =>  inp_feat(11), I3 =>  inp_feat(233), I4 =>  inp_feat(422), I5 =>  inp_feat(501), I6 =>  inp_feat(483), I7 =>  inp_feat(372)); 
C_11_S_4_L_6_inst : LUT8 generic map(INIT => "1111111110111111110100011111110111001100100000001100110000000000101010101110101011101010111010001110111010100000111011101100000000000000000000100000000000000000000000000000000000000000000000001010000000000000000010000000000000000100000000000100010001000100") port map( O =>C_11_S_4_L_6_out, I0 =>  inp_feat(232), I1 =>  inp_feat(327), I2 =>  inp_feat(6), I3 =>  inp_feat(293), I4 =>  inp_feat(290), I5 =>  inp_feat(142), I6 =>  inp_feat(108), I7 =>  inp_feat(489)); 
C_11_S_4_L_7_inst : LUT8 generic map(INIT => "1111110011101100101110000000000011110000111000000000000000000000101110000000000000111000000000000010001000000000000000000000000010110010000000001000000000000000001000100000000000000010000000001010001000000000001000000000000000100010000000000000000000000000") port map( O =>C_11_S_4_L_7_out, I0 =>  inp_feat(396), I1 =>  inp_feat(288), I2 =>  inp_feat(501), I3 =>  inp_feat(437), I4 =>  inp_feat(398), I5 =>  inp_feat(397), I6 =>  inp_feat(14), I7 =>  inp_feat(199)); 
C_12_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_1_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_2_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_3_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_12_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000000110000000000000011000000000000000000000000000000") port map( O =>C_12_S_4_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(1), I2 =>  inp_feat(147), I3 =>  inp_feat(314), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_0_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_0_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_1_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_1_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_2_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_2_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_3_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_0_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_1_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_2_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_3_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_4_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_5_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_6_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_13_S_4_L_7_inst : LUT8 generic map(INIT => "1111101011001010010000101100000000001010110000000000111111001000100010001000000000000000000000000000000000000000000011110000000011001000110010000100000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_13_S_4_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(36), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_0_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_1_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_2_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_3_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_4_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_5_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_6_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_0_L_7_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_0_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_1_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_2_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_3_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_4_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_5_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_6_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_1_L_7_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_0_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_1_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_2_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_3_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_4_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_5_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_6_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_2_L_7_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_0_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_1_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_2_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_3_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_4_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_5_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_6_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_3_L_7_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_0_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_1_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_2_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_3_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_4_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_5_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_6_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_14_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000010110000000000000000000000000000000000000000000000000000110000000000000000000000000000001010000000000000001000000000000010100000100000000000000000000000") port map( O =>C_14_S_4_L_7_out, I0 =>  inp_feat(264), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(318), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_0_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_1_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_2_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_3_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_15_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100000000000100010000000000010001000000000000000000000000000") port map( O =>C_15_S_4_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(1), I2 =>  inp_feat(0), I3 =>  inp_feat(342), I4 =>  inp_feat(143), I5 =>  inp_feat(199), I6 =>  inp_feat(326), I7 =>  inp_feat(352)); 
C_16_S_0_L_0_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_1_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_2_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_3_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_4_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_5_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_6_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_0_L_7_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_0_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_1_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_2_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_3_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_4_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_5_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_6_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_1_L_7_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_1_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_0_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_1_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_2_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_3_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_4_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_5_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_6_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_2_L_7_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_2_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_0_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_1_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_2_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_3_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_4_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_5_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_6_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_3_L_7_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_3_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_0_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_1_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_2_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_3_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_4_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_5_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_6_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_16_S_4_L_7_inst : LUT8 generic map(INIT => "1110111010000010101011100000101011001101000000001000100000000000110111110000001011101110000010101110001100001000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_16_S_4_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(136), I2 =>  inp_feat(448), I3 =>  inp_feat(389), I4 =>  inp_feat(90), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_0_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_1_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_2_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_3_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_0_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_1_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_2_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_3_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_4_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_6_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_17_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000100010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100010000000000000000000") port map( O =>C_17_S_4_L_7_out, I0 =>  inp_feat(2), I1 =>  inp_feat(176), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_18_S_0_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_0_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_18_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111110100111100001000000001110100010101000000000000000000111111101111100000000000000000001100000001000000100000000000000011001000001000000000000000000000000000001011000100000000000000001110110011110000100000000000000011010000111101001000000000000000") port map( O =>C_18_S_0_L_1_out, I0 =>  inp_feat(448), I1 =>  inp_feat(259), I2 =>  inp_feat(262), I3 =>  inp_feat(467), I4 =>  inp_feat(287), I5 =>  inp_feat(78), I6 =>  inp_feat(176), I7 =>  inp_feat(475)); 
C_18_S_0_L_2_inst : LUT8 generic map(INIT => "1000000011000000111000101100000011111110110100001101110000000000111010001010000011000100000000001010000010110000100001000000000010101000100000001010110010100000111100001111000010111100100000001100100000000000100011000000000010101000000000001010100000000000") port map( O =>C_18_S_0_L_2_out, I0 =>  inp_feat(227), I1 =>  inp_feat(473), I2 =>  inp_feat(162), I3 =>  inp_feat(307), I4 =>  inp_feat(228), I5 =>  inp_feat(364), I6 =>  inp_feat(180), I7 =>  inp_feat(472)); 
C_18_S_0_L_3_inst : LUT8 generic map(INIT => "1111110011111110110010001100110011110100111101000000000000000000100010000000000000000000000000001010000000000000000000000000000011000000100000001000100000000000110100000000000001010000000000001000000000000000100000000000000011000000000000000000000000000000") port map( O =>C_18_S_0_L_3_out, I0 =>  inp_feat(493), I1 =>  inp_feat(213), I2 =>  inp_feat(78), I3 =>  inp_feat(484), I4 =>  inp_feat(230), I5 =>  inp_feat(372), I6 =>  inp_feat(16), I7 =>  inp_feat(205)); 
C_18_S_0_L_4_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_18_S_0_L_4_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_18_S_0_L_5_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_18_S_0_L_5_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_18_S_0_L_6_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_18_S_0_L_6_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_18_S_0_L_7_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_18_S_0_L_7_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_18_S_1_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_1_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_18_S_1_L_1_inst : LUT8 generic map(INIT => "1111101110111010110010000001100011111010101010100100100000000000111000000000000001010000000000000000000000000000000000000000000011111010000010000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_1_L_1_out, I0 =>  inp_feat(307), I1 =>  inp_feat(358), I2 =>  inp_feat(283), I3 =>  inp_feat(78), I4 =>  inp_feat(271), I5 =>  inp_feat(270), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_18_S_1_L_2_inst : LUT8 generic map(INIT => "1000100011001000110011001010000010001000100000001100110000000000101010101010000010101111101000101000100011000000000000000000000000001010110010001010000010100000100010000000000000000000000000000010100010000000001000001000000000001000000000000000000000000000") port map( O =>C_18_S_1_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(113), I3 =>  inp_feat(224), I4 =>  inp_feat(221), I5 =>  inp_feat(345), I6 =>  inp_feat(4), I7 =>  inp_feat(273)); 
C_18_S_1_L_3_inst : LUT8 generic map(INIT => "1110110010101100111011001010000011101100101011000000100000000000000001000010000011101100101000000010000000100000000000000000000010000000100010001100100010001000100000001000110010000000100010000000000000000000100000001000000000000000000000001000000000000000") port map( O =>C_18_S_1_L_3_out, I0 =>  inp_feat(466), I1 =>  inp_feat(363), I2 =>  inp_feat(427), I3 =>  inp_feat(467), I4 =>  inp_feat(289), I5 =>  inp_feat(324), I6 =>  inp_feat(500), I7 =>  inp_feat(455)); 
C_18_S_1_L_4_inst : LUT8 generic map(INIT => "1111110111111101111001001100010011000100110011001010110011001100111101011111100010100000100000001010000010101000000000000000000001010101110101011100000011000000000000000000000000100000000000001000000011000000111000001110000000000000000000000000000000000000") port map( O =>C_18_S_1_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(195), I2 =>  inp_feat(205), I3 =>  inp_feat(41), I4 =>  inp_feat(259), I5 =>  inp_feat(34), I6 =>  inp_feat(336), I7 =>  inp_feat(162)); 
C_18_S_1_L_5_inst : LUT8 generic map(INIT => "1111111011111011100111111001000000111111100000001101111100000000111110101111001010010000100000001011000110000000110100001000000001101110111111111000100000000000000000000000000000000000000000001010101010100010100000000000000000000000000000000000000000000000") port map( O =>C_18_S_1_L_5_out, I0 =>  inp_feat(362), I1 =>  inp_feat(81), I2 =>  inp_feat(260), I3 =>  inp_feat(107), I4 =>  inp_feat(215), I5 =>  inp_feat(363), I6 =>  inp_feat(56), I7 =>  inp_feat(457)); 
C_18_S_1_L_6_inst : LUT8 generic map(INIT => "1111101111110000111010100010000011111110101100001010101000100000101010000010000000100000000000000000000000000000000000000000000011000000000000000100100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_1_L_6_out, I0 =>  inp_feat(25), I1 =>  inp_feat(228), I2 =>  inp_feat(3), I3 =>  inp_feat(20), I4 =>  inp_feat(40), I5 =>  inp_feat(425), I6 =>  inp_feat(271), I7 =>  inp_feat(101)); 
C_18_S_1_L_7_inst : LUT8 generic map(INIT => "1111011111100000111101111110000001000000110000001110000011000000111100101010000010110000101000000010000000000000101000001010000010100000101000001000000010100000000000000000000000000000000000000000000010100000001000000000000000000000100000000000000000000000") port map( O =>C_18_S_1_L_7_out, I0 =>  inp_feat(395), I1 =>  inp_feat(472), I2 =>  inp_feat(389), I3 =>  inp_feat(229), I4 =>  inp_feat(228), I5 =>  inp_feat(367), I6 =>  inp_feat(226), I7 =>  inp_feat(307)); 
C_18_S_2_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_2_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_18_S_2_L_1_inst : LUT8 generic map(INIT => "1111101110111010110010000001100011111010101010100100100000000000111000000000000001010000000000000000000000000000000000000000000011111010000010000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_2_L_1_out, I0 =>  inp_feat(307), I1 =>  inp_feat(358), I2 =>  inp_feat(283), I3 =>  inp_feat(78), I4 =>  inp_feat(271), I5 =>  inp_feat(270), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_18_S_2_L_2_inst : LUT8 generic map(INIT => "1000100011001000110011001010000010001000100000001100110000000000101010101010000010101111101000101000100011000000000000000000000000001010110010001010000010100000100010000000000000000000000000000010100010000000001000001000000000001000000000000000000000000000") port map( O =>C_18_S_2_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(113), I3 =>  inp_feat(224), I4 =>  inp_feat(221), I5 =>  inp_feat(345), I6 =>  inp_feat(4), I7 =>  inp_feat(273)); 
C_18_S_2_L_3_inst : LUT8 generic map(INIT => "1110110010101100111011001010000011101100101011000000100000000000000001000010000011101100101000000010000000100000000000000000000010000000100010001100100010001000100000001000110010000000100010000000000000000000100000001000000000000000000000001000000000000000") port map( O =>C_18_S_2_L_3_out, I0 =>  inp_feat(466), I1 =>  inp_feat(363), I2 =>  inp_feat(427), I3 =>  inp_feat(467), I4 =>  inp_feat(289), I5 =>  inp_feat(324), I6 =>  inp_feat(500), I7 =>  inp_feat(455)); 
C_18_S_2_L_4_inst : LUT8 generic map(INIT => "1111110111111101111001001100010011000100110011001010110011001100111101011111100010100000100000001010000010101000000000000000000001010101110101011100000011000000000000000000000000100000000000001000000011000000111000001110000000000000000000000000000000000000") port map( O =>C_18_S_2_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(195), I2 =>  inp_feat(205), I3 =>  inp_feat(41), I4 =>  inp_feat(259), I5 =>  inp_feat(34), I6 =>  inp_feat(336), I7 =>  inp_feat(162)); 
C_18_S_2_L_5_inst : LUT8 generic map(INIT => "1111111011111011100111111001000000111111100000001101111100000000111110101111001010010000100000001011000110000000110100001000000001101110111111111000100000000000000000000000000000000000000000001010101010100010100000000000000000000000000000000000000000000000") port map( O =>C_18_S_2_L_5_out, I0 =>  inp_feat(362), I1 =>  inp_feat(81), I2 =>  inp_feat(260), I3 =>  inp_feat(107), I4 =>  inp_feat(215), I5 =>  inp_feat(363), I6 =>  inp_feat(56), I7 =>  inp_feat(457)); 
C_18_S_2_L_6_inst : LUT8 generic map(INIT => "1110001011101010101000001010101010101010000000001000000010000000110010001100100000000000000000000000000000000000000000000000000011100010001000101110000000100010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_2_L_6_out, I0 =>  inp_feat(188), I1 =>  inp_feat(79), I2 =>  inp_feat(98), I3 =>  inp_feat(224), I4 =>  inp_feat(40), I5 =>  inp_feat(425), I6 =>  inp_feat(271), I7 =>  inp_feat(101)); 
C_18_S_2_L_7_inst : LUT8 generic map(INIT => "1100100011101000001010001111101010101010101010001000000010100000110010001010000010000000111100001010100010100000000000000000000000001001101010000000000011101010101110101010101000000000000010001100000010101000110000001100100010000000101010100000000000000000") port map( O =>C_18_S_2_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(40), I2 =>  inp_feat(356), I3 =>  inp_feat(221), I4 =>  inp_feat(237), I5 =>  inp_feat(358), I6 =>  inp_feat(267), I7 =>  inp_feat(285)); 
C_18_S_3_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_3_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_18_S_3_L_1_inst : LUT8 generic map(INIT => "1111101110111010110010000001100011111010101010100100100000000000111000000000000001010000000000000000000000000000000000000000000011111010000010000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_3_L_1_out, I0 =>  inp_feat(307), I1 =>  inp_feat(358), I2 =>  inp_feat(283), I3 =>  inp_feat(78), I4 =>  inp_feat(271), I5 =>  inp_feat(270), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_18_S_3_L_2_inst : LUT8 generic map(INIT => "1000100011001000110011001010000010001000100000001100110000000000101010101010000010101111101000101000100011000000000000000000000000001010110010001010000010100000100010000000000000000000000000000010100010000000001000001000000000001000000000000000000000000000") port map( O =>C_18_S_3_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(113), I3 =>  inp_feat(224), I4 =>  inp_feat(221), I5 =>  inp_feat(345), I6 =>  inp_feat(4), I7 =>  inp_feat(273)); 
C_18_S_3_L_3_inst : LUT8 generic map(INIT => "1011111010100010101010101010101100100010100000001010001010100010111010101010000011001000100000001000000010100000000000000000000000100011101110101110111111111111000000000000000000001010111111110010011010100000000000001111000000000000000000000000000000010000") port map( O =>C_18_S_3_L_3_out, I0 =>  inp_feat(511), I1 =>  inp_feat(212), I2 =>  inp_feat(94), I3 =>  inp_feat(180), I4 =>  inp_feat(289), I5 =>  inp_feat(500), I6 =>  inp_feat(428), I7 =>  inp_feat(455)); 
C_18_S_3_L_4_inst : LUT8 generic map(INIT => "1010101010100010111010001010000010100010101000000010001010000000110010001000000011000000100000000000000000000000000000001000000010100010100000001000100000000000100000001000000000000000100000001000100010000000000000000000000010000000100000000000000010000000") port map( O =>C_18_S_3_L_4_out, I0 =>  inp_feat(63), I1 =>  inp_feat(315), I2 =>  inp_feat(78), I3 =>  inp_feat(95), I4 =>  inp_feat(474), I5 =>  inp_feat(125), I6 =>  inp_feat(483), I7 =>  inp_feat(98)); 
C_18_S_3_L_5_inst : LUT8 generic map(INIT => "1111111100101000010111010000010011111111000000001100111111000000000011101000110010111110000011000000110100000000100011001000010011111010100000001101000000000000101011100000000000001000000000001100110000000000110011000000000000001000000000000000100000000000") port map( O =>C_18_S_3_L_5_out, I0 =>  inp_feat(344), I1 =>  inp_feat(356), I2 =>  inp_feat(221), I3 =>  inp_feat(511), I4 =>  inp_feat(331), I5 =>  inp_feat(293), I6 =>  inp_feat(56), I7 =>  inp_feat(176)); 
C_18_S_3_L_6_inst : LUT8 generic map(INIT => "1111110011110000101110111010000010001000001000000011000010100000101010001010000011101000101000000000000000000000000000000000000010000000100000001000000000000000000000000000000000000000000000001100000010000000110000001000000000000000000000000000000000000000") port map( O =>C_18_S_3_L_6_out, I0 =>  inp_feat(230), I1 =>  inp_feat(171), I2 =>  inp_feat(292), I3 =>  inp_feat(356), I4 =>  inp_feat(4), I5 =>  inp_feat(162), I6 =>  inp_feat(436), I7 =>  inp_feat(213)); 
C_18_S_3_L_7_inst : LUT8 generic map(INIT => "1110101010100010111010000000000010101000101000101100100000100001111011110000000011000000000000001010000000100000011000000000000111001000000000001010100000000000100000000000100000001000001000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_3_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(195), I2 =>  inp_feat(362), I3 =>  inp_feat(57), I4 =>  inp_feat(259), I5 =>  inp_feat(78), I6 =>  inp_feat(455), I7 =>  inp_feat(271)); 
C_18_S_4_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_4_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_18_S_4_L_1_inst : LUT8 generic map(INIT => "1110101011111010101010101010101010110000101110100000000010100010101000000000000000000000000000000000000000000000000000000000000010100000100000000010000010000000101000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_18_S_4_L_1_out, I0 =>  inp_feat(389), I1 =>  inp_feat(107), I2 =>  inp_feat(511), I3 =>  inp_feat(245), I4 =>  inp_feat(367), I5 =>  inp_feat(195), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_18_S_4_L_2_inst : LUT8 generic map(INIT => "1111000011010000000001000000000011001100110111000000000000000000110000001101000000000000000000001000110001010100000000000000000011100000111000001100110010000000110011001100110011001100000000000000000000000000000010000000000010001000110001000000100000000000") port map( O =>C_18_S_4_L_2_out, I0 =>  inp_feat(493), I1 =>  inp_feat(24), I2 =>  inp_feat(475), I3 =>  inp_feat(195), I4 =>  inp_feat(371), I5 =>  inp_feat(176), I6 =>  inp_feat(78), I7 =>  inp_feat(4)); 
C_18_S_4_L_3_inst : LUT8 generic map(INIT => "1111111111001010111011001100000010100000000000001010000000000000111011001110100010100000100000001010000010100000101000000000000011000000100000000100000010000000000000000000000000000000000000001000000011000000000000001000000010000000100000000000000000000000") port map( O =>C_18_S_4_L_3_out, I0 =>  inp_feat(287), I1 =>  inp_feat(24), I2 =>  inp_feat(195), I3 =>  inp_feat(78), I4 =>  inp_feat(345), I5 =>  inp_feat(20), I6 =>  inp_feat(228), I7 =>  inp_feat(510)); 
C_18_S_4_L_4_inst : LUT8 generic map(INIT => "1110000011001100101010001010100011001000100011001100100000000000110000001100000000000000000000000000000000000000000000000000000011101000000000001000000000000000111000000000000011100000000000001100010000000000000000000000000001010001000000000000000000000000") port map( O =>C_18_S_4_L_4_out, I0 =>  inp_feat(134), I1 =>  inp_feat(162), I2 =>  inp_feat(511), I3 =>  inp_feat(456), I4 =>  inp_feat(5), I5 =>  inp_feat(455), I6 =>  inp_feat(3), I7 =>  inp_feat(427)); 
C_18_S_4_L_5_inst : LUT8 generic map(INIT => "1111111111101111111100010101000011111101000000001111000100000000111011100000111010000000000000001100110000000100000000000000000010000000010000001101000001110101000000000000000010000000000000001000000000000000100000001011011000000000000000000000000000000000") port map( O =>C_18_S_4_L_5_out, I0 =>  inp_feat(212), I1 =>  inp_feat(6), I2 =>  inp_feat(367), I3 =>  inp_feat(78), I4 =>  inp_feat(427), I5 =>  inp_feat(205), I6 =>  inp_feat(259), I7 =>  inp_feat(136)); 
C_18_S_4_L_6_inst : LUT8 generic map(INIT => "1111101011111000111110001101000010101000100010000000100000000000111110001101000000000000000000001010000010000000000000000000000010100000000000000011100000000000101010000000000010001000000000001011000000000000001000000000000010100000000000000010000000000000") port map( O =>C_18_S_4_L_6_out, I0 =>  inp_feat(367), I1 =>  inp_feat(78), I2 =>  inp_feat(213), I3 =>  inp_feat(154), I4 =>  inp_feat(286), I5 =>  inp_feat(359), I6 =>  inp_feat(245), I7 =>  inp_feat(98)); 
C_18_S_4_L_7_inst : LUT8 generic map(INIT => "1111111111001101101010101000000011001000110000001000000000000000111010001000000010111000000000001100000000000000000000000000000011101010000000001000000000000000111010101100000010000000000000001010000000000000100000000000000011000000110000001000000000000000") port map( O =>C_18_S_4_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(78), I2 =>  inp_feat(151), I3 =>  inp_feat(205), I4 =>  inp_feat(356), I5 =>  inp_feat(234), I6 =>  inp_feat(307), I7 =>  inp_feat(82)); 
C_19_S_0_L_0_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_0_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_1_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_1_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_2_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_2_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_3_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_3_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_4_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_4_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_5_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_5_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_6_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_6_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_0_L_7_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_0_L_7_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_0_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_0_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_1_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_1_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_2_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_2_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_3_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_3_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_4_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_4_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_5_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_5_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_6_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_6_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_1_L_7_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_1_L_7_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_0_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_0_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_1_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_1_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_2_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_2_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_3_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_3_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_4_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_4_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_5_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_5_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_6_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_6_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_2_L_7_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_2_L_7_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_0_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_0_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_1_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_1_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_2_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_2_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_3_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_3_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_4_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_4_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_5_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_5_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_6_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_6_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_3_L_7_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_3_L_7_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_0_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_0_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_1_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_1_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_2_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_2_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_3_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_3_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_4_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_4_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_5_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_5_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_6_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_6_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_19_S_4_L_7_inst : LUT8 generic map(INIT => "1111110101110101111110011011010110100000001000101010000000100000111010101010000011101010101010100000000000000000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_19_S_4_L_7_out, I0 =>  inp_feat(28), I1 =>  inp_feat(228), I2 =>  inp_feat(98), I3 =>  inp_feat(78), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_20_S_0_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_20_S_0_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_20_S_0_L_1_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_1_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_0_L_2_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_0_L_3_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_3_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_0_L_4_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_4_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_0_L_5_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_5_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_0_L_6_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_6_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_0_L_7_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_0_L_7_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_20_S_1_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_20_S_1_L_1_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_1_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_2_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_3_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_3_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_4_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_4_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_5_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_5_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_6_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_6_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_1_L_7_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_20_S_1_L_7_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_20_S_2_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_20_S_2_L_1_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_1_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_2_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_2_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_3_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_4_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_5_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_6_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_6_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_2_L_7_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_2_L_7_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_20_S_3_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_20_S_3_L_1_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_1_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_2_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_2_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_3_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_4_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_5_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_6_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_6_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_3_L_7_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_3_L_7_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_20_S_4_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_20_S_4_L_1_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_1_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_2_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_2_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_3_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_4_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_5_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_6_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_6_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_20_S_4_L_7_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_20_S_4_L_7_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_21_S_0_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_0_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_21_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111110100111100001000000001110100010101000000000000000000111111101111100000000000000000001100000001000000100000000000000011001000001000000000000000000000000000001011000100000000000000001110110011110000100000000000000011010000111101001000000000000000") port map( O =>C_21_S_0_L_1_out, I0 =>  inp_feat(448), I1 =>  inp_feat(259), I2 =>  inp_feat(262), I3 =>  inp_feat(467), I4 =>  inp_feat(287), I5 =>  inp_feat(78), I6 =>  inp_feat(176), I7 =>  inp_feat(475)); 
C_21_S_0_L_2_inst : LUT8 generic map(INIT => "1000000011000000111000101100000011111110110100001101110000000000111010001010000011000100000000001010000010110000100001000000000010101000100000001010110010100000111100001111000010111100100000001100100000000000100011000000000010101000000000001010100000000000") port map( O =>C_21_S_0_L_2_out, I0 =>  inp_feat(227), I1 =>  inp_feat(473), I2 =>  inp_feat(162), I3 =>  inp_feat(307), I4 =>  inp_feat(228), I5 =>  inp_feat(364), I6 =>  inp_feat(180), I7 =>  inp_feat(472)); 
C_21_S_0_L_3_inst : LUT8 generic map(INIT => "1111110011111110110010001100110011110100111101000000000000000000100010000000000000000000000000001010000000000000000000000000000011000000100000001000100000000000110100000000000001010000000000001000000000000000100000000000000011000000000000000000000000000000") port map( O =>C_21_S_0_L_3_out, I0 =>  inp_feat(493), I1 =>  inp_feat(213), I2 =>  inp_feat(78), I3 =>  inp_feat(484), I4 =>  inp_feat(230), I5 =>  inp_feat(372), I6 =>  inp_feat(16), I7 =>  inp_feat(205)); 
C_21_S_0_L_4_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_21_S_0_L_4_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_21_S_0_L_5_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_21_S_0_L_5_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_21_S_0_L_6_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_21_S_0_L_6_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_21_S_0_L_7_inst : LUT8 generic map(INIT => "1111100011101000111110000100000011111000110010001101100000000000000100000000000001110000001000001100000000000000111110000000000000100000000000001111000000000000000010000000000001001000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_21_S_0_L_7_out, I0 =>  inp_feat(171), I1 =>  inp_feat(473), I2 =>  inp_feat(213), I3 =>  inp_feat(117), I4 =>  inp_feat(38), I5 =>  inp_feat(387), I6 =>  inp_feat(511), I7 =>  inp_feat(510)); 
C_21_S_1_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_1_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_21_S_1_L_1_inst : LUT8 generic map(INIT => "1111101110111010110010000001100011111010101010100100100000000000111000000000000001010000000000000000000000000000000000000000000011111010000010000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_1_L_1_out, I0 =>  inp_feat(307), I1 =>  inp_feat(358), I2 =>  inp_feat(283), I3 =>  inp_feat(78), I4 =>  inp_feat(271), I5 =>  inp_feat(270), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_21_S_1_L_2_inst : LUT8 generic map(INIT => "1000100011001000110011001010000010001000100000001100110000000000101010101010000010101111101000101000100011000000000000000000000000001010110010001010000010100000100010000000000000000000000000000010100010000000001000001000000000001000000000000000000000000000") port map( O =>C_21_S_1_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(113), I3 =>  inp_feat(224), I4 =>  inp_feat(221), I5 =>  inp_feat(345), I6 =>  inp_feat(4), I7 =>  inp_feat(273)); 
C_21_S_1_L_3_inst : LUT8 generic map(INIT => "1110110010101100111011001010000011101100101011000000100000000000000001000010000011101100101000000010000000100000000000000000000010000000100010001100100010001000100000001000110010000000100010000000000000000000100000001000000000000000000000001000000000000000") port map( O =>C_21_S_1_L_3_out, I0 =>  inp_feat(466), I1 =>  inp_feat(363), I2 =>  inp_feat(427), I3 =>  inp_feat(467), I4 =>  inp_feat(289), I5 =>  inp_feat(324), I6 =>  inp_feat(500), I7 =>  inp_feat(455)); 
C_21_S_1_L_4_inst : LUT8 generic map(INIT => "1111110111111101111001001100010011000100110011001010110011001100111101011111100010100000100000001010000010101000000000000000000001010101110101011100000011000000000000000000000000100000000000001000000011000000111000001110000000000000000000000000000000000000") port map( O =>C_21_S_1_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(195), I2 =>  inp_feat(205), I3 =>  inp_feat(41), I4 =>  inp_feat(259), I5 =>  inp_feat(34), I6 =>  inp_feat(336), I7 =>  inp_feat(162)); 
C_21_S_1_L_5_inst : LUT8 generic map(INIT => "1111111011111011100111111001000000111111100000001101111100000000111110101111001010010000100000001011000110000000110100001000000001101110111111111000100000000000000000000000000000000000000000001010101010100010100000000000000000000000000000000000000000000000") port map( O =>C_21_S_1_L_5_out, I0 =>  inp_feat(362), I1 =>  inp_feat(81), I2 =>  inp_feat(260), I3 =>  inp_feat(107), I4 =>  inp_feat(215), I5 =>  inp_feat(363), I6 =>  inp_feat(56), I7 =>  inp_feat(457)); 
C_21_S_1_L_6_inst : LUT8 generic map(INIT => "1111101111110000111010100010000011111110101100001010101000100000101010000010000000100000000000000000000000000000000000000000000011000000000000000100100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_1_L_6_out, I0 =>  inp_feat(25), I1 =>  inp_feat(228), I2 =>  inp_feat(3), I3 =>  inp_feat(20), I4 =>  inp_feat(40), I5 =>  inp_feat(425), I6 =>  inp_feat(271), I7 =>  inp_feat(101)); 
C_21_S_1_L_7_inst : LUT8 generic map(INIT => "1111011111100000111101111110000001000000110000001110000011000000111100101010000010110000101000000010000000000000101000001010000010100000101000001000000010100000000000000000000000000000000000000000000010100000001000000000000000000000100000000000000000000000") port map( O =>C_21_S_1_L_7_out, I0 =>  inp_feat(395), I1 =>  inp_feat(472), I2 =>  inp_feat(389), I3 =>  inp_feat(229), I4 =>  inp_feat(228), I5 =>  inp_feat(367), I6 =>  inp_feat(226), I7 =>  inp_feat(307)); 
C_21_S_2_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_2_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_21_S_2_L_1_inst : LUT8 generic map(INIT => "1111101110111010110010000001100011111010101010100100100000000000111000000000000001010000000000000000000000000000000000000000000011111010000010000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_2_L_1_out, I0 =>  inp_feat(307), I1 =>  inp_feat(358), I2 =>  inp_feat(283), I3 =>  inp_feat(78), I4 =>  inp_feat(271), I5 =>  inp_feat(270), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_21_S_2_L_2_inst : LUT8 generic map(INIT => "1000100011001000110011001010000010001000100000001100110000000000101010101010000010101111101000101000100011000000000000000000000000001010110010001010000010100000100010000000000000000000000000000010100010000000001000001000000000001000000000000000000000000000") port map( O =>C_21_S_2_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(113), I3 =>  inp_feat(224), I4 =>  inp_feat(221), I5 =>  inp_feat(345), I6 =>  inp_feat(4), I7 =>  inp_feat(273)); 
C_21_S_2_L_3_inst : LUT8 generic map(INIT => "1110110010101100111011001010000011101100101011000000100000000000000001000010000011101100101000000010000000100000000000000000000010000000100010001100100010001000100000001000110010000000100010000000000000000000100000001000000000000000000000001000000000000000") port map( O =>C_21_S_2_L_3_out, I0 =>  inp_feat(466), I1 =>  inp_feat(363), I2 =>  inp_feat(427), I3 =>  inp_feat(467), I4 =>  inp_feat(289), I5 =>  inp_feat(324), I6 =>  inp_feat(500), I7 =>  inp_feat(455)); 
C_21_S_2_L_4_inst : LUT8 generic map(INIT => "1111110111111101111001001100010011000100110011001010110011001100111101011111100010100000100000001010000010101000000000000000000001010101110101011100000011000000000000000000000000100000000000001000000011000000111000001110000000000000000000000000000000000000") port map( O =>C_21_S_2_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(195), I2 =>  inp_feat(205), I3 =>  inp_feat(41), I4 =>  inp_feat(259), I5 =>  inp_feat(34), I6 =>  inp_feat(336), I7 =>  inp_feat(162)); 
C_21_S_2_L_5_inst : LUT8 generic map(INIT => "1111111011111011100111111001000000111111100000001101111100000000111110101111001010010000100000001011000110000000110100001000000001101110111111111000100000000000000000000000000000000000000000001010101010100010100000000000000000000000000000000000000000000000") port map( O =>C_21_S_2_L_5_out, I0 =>  inp_feat(362), I1 =>  inp_feat(81), I2 =>  inp_feat(260), I3 =>  inp_feat(107), I4 =>  inp_feat(215), I5 =>  inp_feat(363), I6 =>  inp_feat(56), I7 =>  inp_feat(457)); 
C_21_S_2_L_6_inst : LUT8 generic map(INIT => "1110001011101010101000001010101010101010000000001000000010000000110010001100100000000000000000000000000000000000000000000000000011100010001000101110000000100010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_2_L_6_out, I0 =>  inp_feat(188), I1 =>  inp_feat(79), I2 =>  inp_feat(98), I3 =>  inp_feat(224), I4 =>  inp_feat(40), I5 =>  inp_feat(425), I6 =>  inp_feat(271), I7 =>  inp_feat(101)); 
C_21_S_2_L_7_inst : LUT8 generic map(INIT => "1100100011101000001010001111101010101010101010001000000010100000110010001010000010000000111100001010100010100000000000000000000000001001101010000000000011101010101110101010101000000000000010001100000010101000110000001100100010000000101010100000000000000000") port map( O =>C_21_S_2_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(40), I2 =>  inp_feat(356), I3 =>  inp_feat(221), I4 =>  inp_feat(237), I5 =>  inp_feat(358), I6 =>  inp_feat(267), I7 =>  inp_feat(285)); 
C_21_S_3_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_3_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_21_S_3_L_1_inst : LUT8 generic map(INIT => "1111101110111010110010000001100011111010101010100100100000000000111000000000000001010000000000000000000000000000000000000000000011111010000010000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_3_L_1_out, I0 =>  inp_feat(307), I1 =>  inp_feat(358), I2 =>  inp_feat(283), I3 =>  inp_feat(78), I4 =>  inp_feat(271), I5 =>  inp_feat(270), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_21_S_3_L_2_inst : LUT8 generic map(INIT => "1000100011001000110011001010000010001000100000001100110000000000101010101010000010101111101000101000100011000000000000000000000000001010110010001010000010100000100010000000000000000000000000000010100010000000001000001000000000001000000000000000000000000000") port map( O =>C_21_S_3_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(113), I3 =>  inp_feat(224), I4 =>  inp_feat(221), I5 =>  inp_feat(345), I6 =>  inp_feat(4), I7 =>  inp_feat(273)); 
C_21_S_3_L_3_inst : LUT8 generic map(INIT => "1011111010100010101010101010101100100010100000001010001010100010111010101010000011001000100000001000000010100000000000000000000000100011101110101110111111111111000000000000000000001010111111110010011010100000000000001111000000000000000000000000000000010000") port map( O =>C_21_S_3_L_3_out, I0 =>  inp_feat(511), I1 =>  inp_feat(212), I2 =>  inp_feat(94), I3 =>  inp_feat(180), I4 =>  inp_feat(289), I5 =>  inp_feat(500), I6 =>  inp_feat(428), I7 =>  inp_feat(455)); 
C_21_S_3_L_4_inst : LUT8 generic map(INIT => "1010101010100010111010001010000010100010101000000010001010000000110010001000000011000000100000000000000000000000000000001000000010100010100000001000100000000000100000001000000000000000100000001000100010000000000000000000000010000000100000000000000010000000") port map( O =>C_21_S_3_L_4_out, I0 =>  inp_feat(63), I1 =>  inp_feat(315), I2 =>  inp_feat(78), I3 =>  inp_feat(95), I4 =>  inp_feat(474), I5 =>  inp_feat(125), I6 =>  inp_feat(483), I7 =>  inp_feat(98)); 
C_21_S_3_L_5_inst : LUT8 generic map(INIT => "1111111100101000010111010000010011111111000000001100111111000000000011101000110010111110000011000000110100000000100011001000010011111010100000001101000000000000101011100000000000001000000000001100110000000000110011000000000000001000000000000000100000000000") port map( O =>C_21_S_3_L_5_out, I0 =>  inp_feat(344), I1 =>  inp_feat(356), I2 =>  inp_feat(221), I3 =>  inp_feat(511), I4 =>  inp_feat(331), I5 =>  inp_feat(293), I6 =>  inp_feat(56), I7 =>  inp_feat(176)); 
C_21_S_3_L_6_inst : LUT8 generic map(INIT => "1111110011110000101110111010000010001000001000000011000010100000101010001010000011101000101000000000000000000000000000000000000010000000100000001000000000000000000000000000000000000000000000001100000010000000110000001000000000000000000000000000000000000000") port map( O =>C_21_S_3_L_6_out, I0 =>  inp_feat(230), I1 =>  inp_feat(171), I2 =>  inp_feat(292), I3 =>  inp_feat(356), I4 =>  inp_feat(4), I5 =>  inp_feat(162), I6 =>  inp_feat(436), I7 =>  inp_feat(213)); 
C_21_S_3_L_7_inst : LUT8 generic map(INIT => "1110101010100010111010000000000010101000101000101100100000100001111011110000000011000000000000001010000000100000011000000000000111001000000000001010100000000000100000000000100000001000001000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_3_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(195), I2 =>  inp_feat(362), I3 =>  inp_feat(57), I4 =>  inp_feat(259), I5 =>  inp_feat(78), I6 =>  inp_feat(455), I7 =>  inp_feat(271)); 
C_21_S_4_L_0_inst : LUT8 generic map(INIT => "1110110001001000101010101000100010001000100010001000100010001000110011100000000011001010100010000000000000000000100010000000100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_4_L_0_out, I0 =>  inp_feat(213), I1 =>  inp_feat(389), I2 =>  inp_feat(107), I3 =>  inp_feat(511), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_21_S_4_L_1_inst : LUT8 generic map(INIT => "1110101011111010101010101010101010110000101110100000000010100010101000000000000000000000000000000000000000000000000000000000000010100000100000000010000010000000101000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_21_S_4_L_1_out, I0 =>  inp_feat(389), I1 =>  inp_feat(107), I2 =>  inp_feat(511), I3 =>  inp_feat(245), I4 =>  inp_feat(367), I5 =>  inp_feat(195), I6 =>  inp_feat(63), I7 =>  inp_feat(16)); 
C_21_S_4_L_2_inst : LUT8 generic map(INIT => "1111000011010000000001000000000011001100110111000000000000000000110000001101000000000000000000001000110001010100000000000000000011100000111000001100110010000000110011001100110011001100000000000000000000000000000010000000000010001000110001000000100000000000") port map( O =>C_21_S_4_L_2_out, I0 =>  inp_feat(493), I1 =>  inp_feat(24), I2 =>  inp_feat(475), I3 =>  inp_feat(195), I4 =>  inp_feat(371), I5 =>  inp_feat(176), I6 =>  inp_feat(78), I7 =>  inp_feat(4)); 
C_21_S_4_L_3_inst : LUT8 generic map(INIT => "1111111111001010111011001100000010100000000000001010000000000000111011001110100010100000100000001010000010100000101000000000000011000000100000000100000010000000000000000000000000000000000000001000000011000000000000001000000010000000100000000000000000000000") port map( O =>C_21_S_4_L_3_out, I0 =>  inp_feat(287), I1 =>  inp_feat(24), I2 =>  inp_feat(195), I3 =>  inp_feat(78), I4 =>  inp_feat(345), I5 =>  inp_feat(20), I6 =>  inp_feat(228), I7 =>  inp_feat(510)); 
C_21_S_4_L_4_inst : LUT8 generic map(INIT => "1110000011001100101010001010100011001000100011001100100000000000110000001100000000000000000000000000000000000000000000000000000011101000000000001000000000000000111000000000000011100000000000001100010000000000000000000000000001010001000000000000000000000000") port map( O =>C_21_S_4_L_4_out, I0 =>  inp_feat(134), I1 =>  inp_feat(162), I2 =>  inp_feat(511), I3 =>  inp_feat(456), I4 =>  inp_feat(5), I5 =>  inp_feat(455), I6 =>  inp_feat(3), I7 =>  inp_feat(427)); 
C_21_S_4_L_5_inst : LUT8 generic map(INIT => "1111111111101111111100010101000011111101000000001111000100000000111011100000111010000000000000001100110000000100000000000000000010000000010000001101000001110101000000000000000010000000000000001000000000000000100000001011011000000000000000000000000000000000") port map( O =>C_21_S_4_L_5_out, I0 =>  inp_feat(212), I1 =>  inp_feat(6), I2 =>  inp_feat(367), I3 =>  inp_feat(78), I4 =>  inp_feat(427), I5 =>  inp_feat(205), I6 =>  inp_feat(259), I7 =>  inp_feat(136)); 
C_21_S_4_L_6_inst : LUT8 generic map(INIT => "1111101011111000111110001101000010101000100010000000100000000000111110001101000000000000000000001010000010000000000000000000000010100000000000000011100000000000101010000000000010001000000000001011000000000000001000000000000010100000000000000010000000000000") port map( O =>C_21_S_4_L_6_out, I0 =>  inp_feat(367), I1 =>  inp_feat(78), I2 =>  inp_feat(213), I3 =>  inp_feat(154), I4 =>  inp_feat(286), I5 =>  inp_feat(359), I6 =>  inp_feat(245), I7 =>  inp_feat(98)); 
C_21_S_4_L_7_inst : LUT8 generic map(INIT => "1111111111001101101010101000000011001000110000001000000000000000111010001000000010111000000000001100000000000000000000000000000011101010000000001000000000000000111010101100000010000000000000001010000000000000100000000000000011000000110000001000000000000000") port map( O =>C_21_S_4_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(78), I2 =>  inp_feat(151), I3 =>  inp_feat(205), I4 =>  inp_feat(356), I5 =>  inp_feat(234), I6 =>  inp_feat(307), I7 =>  inp_feat(82)); 
C_22_S_0_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_22_S_0_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_22_S_0_L_1_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_1_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_0_L_2_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_0_L_3_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_3_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_0_L_4_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_4_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_0_L_5_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_5_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_0_L_6_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_6_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_0_L_7_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_0_L_7_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_22_S_1_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_22_S_1_L_1_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_1_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_2_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_3_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_3_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_4_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_4_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_5_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_5_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_6_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_6_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_1_L_7_inst : LUT8 generic map(INIT => "1110111000101000101011000000000010101110101010100010011000000000111111101010101000101110000000001010101010101010001011100000000001101010000000000000100000010000100011101110110010100000000000001110001000000000001000100001000010100010101100100110001010000000") port map( O =>C_22_S_1_L_7_out, I0 =>  inp_feat(404), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_22_S_2_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_22_S_2_L_1_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_1_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_2_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_2_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_3_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_4_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_5_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_6_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_6_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_2_L_7_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_2_L_7_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_22_S_3_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_22_S_3_L_1_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_1_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_2_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_2_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_3_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_4_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_5_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_6_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_6_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_3_L_7_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_3_L_7_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_0_inst : LUT8 generic map(INIT => "1110111110100010111011101010000011001100000000001100010000000000101111111010001111101111111011100000000000000000110001000100000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_22_S_4_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(293), I2 =>  inp_feat(204), I3 =>  inp_feat(307), I4 =>  inp_feat(245), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_22_S_4_L_1_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_1_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_2_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_2_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_3_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_4_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_5_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_6_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_6_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_22_S_4_L_7_inst : LUT8 generic map(INIT => "1111111100011001101010000000000010001000100010000011101000000000101110001000100010101010000000001011101011001100001010000000000000101000000000000000100000100000001010001010100000100000000000001011100000000000101010000010000000111000111110001010100000010000") port map( O =>C_22_S_4_L_7_out, I0 =>  inp_feat(155), I1 =>  inp_feat(23), I2 =>  inp_feat(221), I3 =>  inp_feat(367), I4 =>  inp_feat(57), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_23_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000110000001000000001000000000000001000000000000000000010000000000000100000111010001110100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000011001000") port map( O =>C_23_S_0_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(228), I2 =>  inp_feat(428), I3 =>  inp_feat(271), I4 =>  inp_feat(511), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_23_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000110000001000000001000000000000001000000000000000000010000000000000100000111010001110100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000011001000") port map( O =>C_23_S_1_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(228), I2 =>  inp_feat(428), I3 =>  inp_feat(271), I4 =>  inp_feat(511), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_23_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_1_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000110000001000000001000000000000001000000000000000000010000000000000100000111010001110100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000011001000") port map( O =>C_23_S_2_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(228), I2 =>  inp_feat(428), I3 =>  inp_feat(271), I4 =>  inp_feat(511), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_23_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000101010100000100000000000000000100000000000000000100000000000000000001010000000000000000000000000000000000000000000000000001010000010001000000000100000001000001000100000000000000000000000100010001010100000000000100010") port map( O =>C_23_S_2_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(40), I2 =>  inp_feat(213), I3 =>  inp_feat(162), I4 =>  inp_feat(29), I5 =>  inp_feat(511), I6 =>  inp_feat(389), I7 =>  inp_feat(134)); 
C_23_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000110000001000000001000000000000001000000000000000000010000000000000100000111010001110100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000011001000") port map( O =>C_23_S_3_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(228), I2 =>  inp_feat(428), I3 =>  inp_feat(271), I4 =>  inp_feat(511), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_23_S_3_L_1_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_1_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_3_L_2_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_2_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_3_L_3_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_3_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_3_L_4_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_4_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_3_L_5_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_5_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_3_L_6_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_6_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_3_L_7_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_3_L_7_out, I0 =>  inp_feat(213), I1 =>  inp_feat(4), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000110000001000000001000000000000001000000000000000000010000000000000100000111010001110100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000011001000") port map( O =>C_23_S_4_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(228), I2 =>  inp_feat(428), I3 =>  inp_feat(271), I4 =>  inp_feat(511), I5 =>  inp_feat(367), I6 =>  inp_feat(195), I7 =>  inp_feat(63)); 
C_23_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000001000000011000000000000000000000000000000010000000000000000001100010001001100000000000000000000000000100000000000000000000000000000000000100000000000000000000000110000000100000000000000000011000000110011000000000000000000") port map( O =>C_23_S_4_L_1_out, I0 =>  inp_feat(213), I1 =>  inp_feat(139), I2 =>  inp_feat(230), I3 =>  inp_feat(234), I4 =>  inp_feat(358), I5 =>  inp_feat(162), I6 =>  inp_feat(136), I7 =>  inp_feat(134)); 
C_23_S_4_L_2_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111100000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_23_S_4_L_2_out, I0 =>  inp_feat(511), I1 =>  inp_feat(509), I2 =>  inp_feat(82), I3 =>  inp_feat(99), I4 =>  inp_feat(322), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_23_S_4_L_3_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111100000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_23_S_4_L_3_out, I0 =>  inp_feat(511), I1 =>  inp_feat(509), I2 =>  inp_feat(82), I3 =>  inp_feat(99), I4 =>  inp_feat(322), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_23_S_4_L_4_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111100000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_23_S_4_L_4_out, I0 =>  inp_feat(511), I1 =>  inp_feat(509), I2 =>  inp_feat(82), I3 =>  inp_feat(99), I4 =>  inp_feat(322), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_23_S_4_L_5_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111100000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_23_S_4_L_5_out, I0 =>  inp_feat(511), I1 =>  inp_feat(509), I2 =>  inp_feat(82), I3 =>  inp_feat(99), I4 =>  inp_feat(322), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_23_S_4_L_6_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111100000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_23_S_4_L_6_out, I0 =>  inp_feat(511), I1 =>  inp_feat(509), I2 =>  inp_feat(82), I3 =>  inp_feat(99), I4 =>  inp_feat(322), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_23_S_4_L_7_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111100000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_23_S_4_L_7_out, I0 =>  inp_feat(511), I1 =>  inp_feat(509), I2 =>  inp_feat(82), I3 =>  inp_feat(99), I4 =>  inp_feat(322), I5 =>  inp_feat(228), I6 =>  inp_feat(176), I7 =>  inp_feat(78)); 
C_24_S_0_L_0_inst : LUT8 generic map(INIT => "1010101111001010111011111100101010111101110011101011101100101010100000001010101010101010101010100010100000100010001010100010101000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_24_S_0_L_0_out, I0 =>  inp_feat(145), I1 =>  inp_feat(62), I2 =>  inp_feat(467), I3 =>  inp_feat(316), I4 =>  inp_feat(413), I5 =>  inp_feat(328), I6 =>  inp_feat(29), I7 =>  inp_feat(299)); 
C_24_S_0_L_1_inst : LUT8 generic map(INIT => "0001110001011101111100001101000011111010101010001111101010011010110000001000000010000000000000001010000000000000100010001000000000011011000000000010000011001100110110100100010111110000110011011100000011001100000000000000110010000000000010001000000000001100") port map( O =>C_24_S_0_L_1_out, I0 =>  inp_feat(290), I1 =>  inp_feat(238), I2 =>  inp_feat(182), I3 =>  inp_feat(416), I4 =>  inp_feat(80), I5 =>  inp_feat(331), I6 =>  inp_feat(148), I7 =>  inp_feat(75)); 
C_24_S_0_L_2_inst : LUT8 generic map(INIT => "0010001011000000101010000010001001100011111001011011100100000000100010001010001010000000000000000000100010000010000000000000000000000000000010101010000000001010011001000000000010100000000000000000000000000000101000000000000010000000000000001010000000000000") port map( O =>C_24_S_0_L_2_out, I0 =>  inp_feat(325), I1 =>  inp_feat(428), I2 =>  inp_feat(509), I3 =>  inp_feat(161), I4 =>  inp_feat(100), I5 =>  inp_feat(220), I6 =>  inp_feat(405), I7 =>  inp_feat(403)); 
C_24_S_0_L_3_inst : LUT8 generic map(INIT => "0111011101110011111000001101010111101101101011110000000001010101100011110010111100110010000100001011111100101011001001000000000011100100111101011010000001010000000010110000000000000000100000001110011101110011011100110001100011111111101111111010110110111110") port map( O =>C_24_S_0_L_3_out, I0 =>  inp_feat(316), I1 =>  inp_feat(290), I2 =>  inp_feat(178), I3 =>  inp_feat(201), I4 =>  inp_feat(308), I5 =>  inp_feat(83), I6 =>  inp_feat(142), I7 =>  inp_feat(373)); 
C_24_S_0_L_4_inst : LUT8 generic map(INIT => "0100010011001111000000000000110011111100000000000000000001001101101111110001000111101100011011110000100000000000000000001111010011011000011101111100000011011101000000000000000000000000011110111100111111010011100100111111011100000000100000000000000011110000") port map( O =>C_24_S_0_L_4_out, I0 =>  inp_feat(290), I1 =>  inp_feat(41), I2 =>  inp_feat(480), I3 =>  inp_feat(488), I4 =>  inp_feat(29), I5 =>  inp_feat(95), I6 =>  inp_feat(105), I7 =>  inp_feat(362)); 
C_24_S_0_L_5_inst : LUT8 generic map(INIT => "1110011000110110111100000001000010111011111111111101100100000000000000000100010000000000000000001000000000000000000000000000000011101100100000000100000000000000101000000000000000000000000000001100000000000000000000000000000010000000000000001000000000000000") port map( O =>C_24_S_0_L_5_out, I0 =>  inp_feat(247), I1 =>  inp_feat(506), I2 =>  inp_feat(29), I3 =>  inp_feat(31), I4 =>  inp_feat(244), I5 =>  inp_feat(7), I6 =>  inp_feat(464), I7 =>  inp_feat(353)); 
C_24_S_0_L_6_inst : LUT8 generic map(INIT => "1100111000001110111011110000001011111110000000001011100010000010010010100000001010101000000000000011011100000010010110100000000011100110000010101110111000000010101001100000001011000010100000100110111000000010011010100000001001101010000000100101001100000010") port map( O =>C_24_S_0_L_6_out, I0 =>  inp_feat(504), I1 =>  inp_feat(15), I2 =>  inp_feat(306), I3 =>  inp_feat(300), I4 =>  inp_feat(265), I5 =>  inp_feat(32), I6 =>  inp_feat(460), I7 =>  inp_feat(290)); 
C_24_S_0_L_7_inst : LUT8 generic map(INIT => "1001110011001000111100001100000011011101110100011111000101010101111110111100000010110001000000001101101101010000011100010100000000100000011110101101000100110011111101000001011111110000000000000011000001110011000100000011001100110011001100110011001100110011") port map( O =>C_24_S_0_L_7_out, I0 =>  inp_feat(420), I1 =>  inp_feat(182), I2 =>  inp_feat(221), I3 =>  inp_feat(290), I4 =>  inp_feat(83), I5 =>  inp_feat(105), I6 =>  inp_feat(353), I7 =>  inp_feat(228)); 
C_24_S_1_L_0_inst : LUT8 generic map(INIT => "1110111111101111001001110010001011001111100011011000111100000100101010110010111100101011001000101011111100001101000000010000000000000100001000100000101000000010100010000000000000001100000000001000100000100010000010000010001010111110000000000000100000000000") port map( O =>C_24_S_1_L_0_out, I0 =>  inp_feat(505), I1 =>  inp_feat(87), I2 =>  inp_feat(478), I3 =>  inp_feat(508), I4 =>  inp_feat(457), I5 =>  inp_feat(200), I6 =>  inp_feat(272), I7 =>  inp_feat(178)); 
C_24_S_1_L_1_inst : LUT8 generic map(INIT => "0111111111111100011111000111110010100000101010000000000010000000111100101111000000000000000000001010000011100000000000000000000010010101100000000100000011000000000000000000000000000000000000001100000011100000110000001100000000000000111000000000000000000000") port map( O =>C_24_S_1_L_1_out, I0 =>  inp_feat(200), I1 =>  inp_feat(100), I2 =>  inp_feat(7), I3 =>  inp_feat(90), I4 =>  inp_feat(211), I5 =>  inp_feat(95), I6 =>  inp_feat(405), I7 =>  inp_feat(178)); 
C_24_S_1_L_2_inst : LUT8 generic map(INIT => "0101101010100000111111010011001011000100000000001001010100010001100011100000100011111111111110110001110010001000111110110000000110000100000010000000101110010011100000000000000000010001000100010000010011011000101111111011011101000000010100011111101111111011") port map( O =>C_24_S_1_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(115), I2 =>  inp_feat(316), I3 =>  inp_feat(259), I4 =>  inp_feat(283), I5 =>  inp_feat(414), I6 =>  inp_feat(420), I7 =>  inp_feat(95)); 
C_24_S_1_L_3_inst : LUT8 generic map(INIT => "1100101011101100101010001000001110101000100001000000100000000000011010001110101100100000001000001111111011011010100000000000000011101010111010001110111011100010111110100101110110101100000000100010000010101111001010100011001111111000011011010100011001101000") port map( O =>C_24_S_1_L_3_out, I0 =>  inp_feat(221), I1 =>  inp_feat(201), I2 =>  inp_feat(373), I3 =>  inp_feat(448), I4 =>  inp_feat(238), I5 =>  inp_feat(187), I6 =>  inp_feat(141), I7 =>  inp_feat(290)); 
C_24_S_1_L_4_inst : LUT8 generic map(INIT => "0110111011111011001010101111001110101110000011110000010000000111100000101001000100110001111111011000100000001111001000000000111100100000101010000010000010000000000010100000111000000000000000000000000000000000001110110010101000000000000010100000000100000010") port map( O =>C_24_S_1_L_4_out, I0 =>  inp_feat(41), I1 =>  inp_feat(316), I2 =>  inp_feat(164), I3 =>  inp_feat(413), I4 =>  inp_feat(210), I5 =>  inp_feat(500), I6 =>  inp_feat(451), I7 =>  inp_feat(144)); 
C_24_S_1_L_5_inst : LUT8 generic map(INIT => "1011111000111000110101001111101000011010010000001101001000000010011100001101101001110010001100100100000001000000010100100010101000001000000000101101101010100010000000000000100000000010001000000000000000000000000100100010101000000000000000000000001010101010") port map( O =>C_24_S_1_L_5_out, I0 =>  inp_feat(331), I1 =>  inp_feat(506), I2 =>  inp_feat(60), I3 =>  inp_feat(40), I4 =>  inp_feat(413), I5 =>  inp_feat(29), I6 =>  inp_feat(322), I7 =>  inp_feat(460)); 
C_24_S_1_L_6_inst : LUT8 generic map(INIT => "0110000111110001101000001011000011110101001000101001010010110000111001000010000010100000111100000101010000100000000000000111000100110000000000010000000010100000000100010000000000000000101100100000000001010000000000001111000000000000001100000000000011110000") port map( O =>C_24_S_1_L_6_out, I0 =>  inp_feat(328), I1 =>  inp_feat(336), I2 =>  inp_feat(179), I3 =>  inp_feat(462), I4 =>  inp_feat(506), I5 =>  inp_feat(493), I6 =>  inp_feat(322), I7 =>  inp_feat(460)); 
C_24_S_1_L_7_inst : LUT8 generic map(INIT => "1100011110001010011101100010001000000000100000100010011110001110000001001010011000010000001000000000011001001100001011110000111010000101100010100000000000000000000010001000100000001000000000000000001100000010000000000000000000000000000000100000000000000000") port map( O =>C_24_S_1_L_7_out, I0 =>  inp_feat(302), I1 =>  inp_feat(452), I2 =>  inp_feat(478), I3 =>  inp_feat(224), I4 =>  inp_feat(180), I5 =>  inp_feat(324), I6 =>  inp_feat(218), I7 =>  inp_feat(120)); 
C_24_S_2_L_0_inst : LUT8 generic map(INIT => "1010101110110101001010011000110111111111110011010000100010010101111101111101000111010101100111111000000100010001000000010001010100000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_24_S_2_L_0_out, I0 =>  inp_feat(61), I1 =>  inp_feat(431), I2 =>  inp_feat(161), I3 =>  inp_feat(200), I4 =>  inp_feat(56), I5 =>  inp_feat(239), I6 =>  inp_feat(194), I7 =>  inp_feat(299)); 
C_24_S_2_L_1_inst : LUT8 generic map(INIT => "1011111011100110111110000010000000100000000000001110000000100000110001000000100010000000000000000000000000000000000000000000000011101110100000101100110011001010001000100010101000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_24_S_2_L_1_out, I0 =>  inp_feat(238), I1 =>  inp_feat(30), I2 =>  inp_feat(340), I3 =>  inp_feat(56), I4 =>  inp_feat(462), I5 =>  inp_feat(18), I6 =>  inp_feat(29), I7 =>  inp_feat(194)); 
C_24_S_2_L_2_inst : LUT8 generic map(INIT => "0111110110100000111010001011000011110101010000000000000000000000110111010000000000001000001000011111010100000000000101010000000011101000101100101110000000110000100010000000000000000000000000001000000000010001000100000000000010001001000000000000000000000000") port map( O =>C_24_S_2_L_2_out, I0 =>  inp_feat(351), I1 =>  inp_feat(302), I2 =>  inp_feat(186), I3 =>  inp_feat(210), I4 =>  inp_feat(405), I5 =>  inp_feat(403), I6 =>  inp_feat(222), I7 =>  inp_feat(247)); 
C_24_S_2_L_3_inst : LUT8 generic map(INIT => "0100100011001000000010001000001001000000000000001000000010001000010110001000000010001000000000000110000010000000000000000000000010001000100000000010101110101010000000001000000000101000001010101010000010000000101100111010101110110000100000001000000000110000") port map( O =>C_24_S_2_L_3_out, I0 =>  inp_feat(277), I1 =>  inp_feat(18), I2 =>  inp_feat(57), I3 =>  inp_feat(173), I4 =>  inp_feat(61), I5 =>  inp_feat(31), I6 =>  inp_feat(385), I7 =>  inp_feat(247)); 
C_24_S_2_L_4_inst : LUT8 generic map(INIT => "1010101100011010100110110000111110101011001100110010111100100111111111110000101010101100000010001100111100000111000010010000101111110001001101001011101100000000100010111110111100001000000000101000110010001000000011000000100000001110000010110000110100001110") port map( O =>C_24_S_2_L_4_out, I0 =>  inp_feat(373), I1 =>  inp_feat(290), I2 =>  inp_feat(5), I3 =>  inp_feat(52), I4 =>  inp_feat(95), I5 =>  inp_feat(367), I6 =>  inp_feat(148), I7 =>  inp_feat(161)); 
C_24_S_2_L_5_inst : LUT8 generic map(INIT => "0011110001111001000000001010000000010000111100100000000000000000101100011111111100000000000000000000000000111000000000000000000011110000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_24_S_2_L_5_out, I0 =>  inp_feat(120), I1 =>  inp_feat(477), I2 =>  inp_feat(42), I3 =>  inp_feat(362), I4 =>  inp_feat(299), I5 =>  inp_feat(467), I6 =>  inp_feat(339), I7 =>  inp_feat(393)); 
C_24_S_2_L_6_inst : LUT8 generic map(INIT => "1101011000110111000010001111111110000011001010111001010111111101100111111101111111111111111111111100111101001111100011110101110101000000010000010000110000000000000000000101000000000000000000000101110101001111111111111111111100000000000000000000000000010000") port map( O =>C_24_S_2_L_6_out, I0 =>  inp_feat(82), I1 =>  inp_feat(52), I2 =>  inp_feat(413), I3 =>  inp_feat(316), I4 =>  inp_feat(161), I5 =>  inp_feat(53), I6 =>  inp_feat(420), I7 =>  inp_feat(144)); 
C_24_S_2_L_7_inst : LUT8 generic map(INIT => "1101111010001100100101110010101111010101000001000101011100001000001000000000000000010000000010001010000000000000000001010000100011100000000000001110000000000000100001000000000001101010000000000000000000000000000000000000000000000000000000000100101000000000") port map( O =>C_24_S_2_L_7_out, I0 =>  inp_feat(161), I1 =>  inp_feat(295), I2 =>  inp_feat(30), I3 =>  inp_feat(393), I4 =>  inp_feat(105), I5 =>  inp_feat(251), I6 =>  inp_feat(300), I7 =>  inp_feat(322)); 
C_24_S_3_L_0_inst : LUT8 generic map(INIT => "1010100000001100011010101001101000001000000011001000100011111100100010100010101000100011000000010000001000001000000000000000000010001000100010100010100111111011000000000000000010001000111111101000001010101010001110111111111100000000000000000000000000000000") port map( O =>C_24_S_3_L_0_out, I0 =>  inp_feat(277), I1 =>  inp_feat(329), I2 =>  inp_feat(480), I3 =>  inp_feat(478), I4 =>  inp_feat(180), I5 =>  inp_feat(256), I6 =>  inp_feat(492), I7 =>  inp_feat(64)); 
C_24_S_3_L_1_inst : LUT8 generic map(INIT => "0010001110001010110001100000000000000010001000100000000000000000111010110010001011000000000000101010000000100010000000000000000011001001001011101100100000000000111001111010001000000000000000001111101010100010111111100000000011110011101010110000000000000010") port map( O =>C_24_S_3_L_1_out, I0 =>  inp_feat(74), I1 =>  inp_feat(135), I2 =>  inp_feat(31), I3 =>  inp_feat(93), I4 =>  inp_feat(18), I5 =>  inp_feat(238), I6 =>  inp_feat(431), I7 =>  inp_feat(478)); 
C_24_S_3_L_2_inst : LUT8 generic map(INIT => "0111111101011110111110000001111000000000000000000001000000000000011110111000001111011111001111110000000000000000000000000000000011010101000000001101010000000100000000000000000000000000000000000000000000000000010101010000010000000000000000000000000000000000") port map( O =>C_24_S_3_L_2_out, I0 =>  inp_feat(362), I1 =>  inp_feat(290), I2 =>  inp_feat(6), I3 =>  inp_feat(43), I4 =>  inp_feat(324), I5 =>  inp_feat(299), I6 =>  inp_feat(467), I7 =>  inp_feat(339)); 
C_24_S_3_L_3_inst : LUT8 generic map(INIT => "0011111011111111001110011100011111100110101100110011000010010001000101111000101100100110000001110010010000000001000010100010000110001111111111110000110110110011101101111011001101101010101100101001111111111111000011110010110101101110101110110000101100110011") port map( O =>C_24_S_3_L_3_out, I0 =>  inp_feat(52), I1 =>  inp_feat(362), I2 =>  inp_feat(382), I3 =>  inp_feat(82), I4 =>  inp_feat(373), I5 =>  inp_feat(500), I6 =>  inp_feat(470), I7 =>  inp_feat(83)); 
C_24_S_3_L_4_inst : LUT8 generic map(INIT => "0111011110110101111011101100100011100000100000001110000000000000111000011111101100000000000000001000000000010000100000000000000000010110000100000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_24_S_3_L_4_out, I0 =>  inp_feat(161), I1 =>  inp_feat(493), I2 =>  inp_feat(262), I3 =>  inp_feat(490), I4 =>  inp_feat(477), I5 =>  inp_feat(393), I6 =>  inp_feat(18), I7 =>  inp_feat(228)); 
C_24_S_3_L_5_inst : LUT8 generic map(INIT => "1100111111011101111110011101110111101110111011001101000000000000010111111101111111010000101101010010001011100000000100000001000001001111110011011000100110001001101110101010000000000001000100000100110001001111000000000001000000000110000000000100000000000001") port map( O =>C_24_S_3_L_5_out, I0 =>  inp_feat(53), I1 =>  inp_feat(467), I2 =>  inp_feat(353), I3 =>  inp_feat(290), I4 =>  inp_feat(239), I5 =>  inp_feat(80), I6 =>  inp_feat(41), I7 =>  inp_feat(339)); 
C_24_S_3_L_6_inst : LUT8 generic map(INIT => "0100100010000011101111101111101110111100100100000000011000000000000000011000001100101100111101100000010000000000000001110011010100001100100010000000110010001000000000000000000000000001000000000000110110000011000011000000111000000111000000010000110000000000") port map( O =>C_24_S_3_L_6_out, I0 =>  inp_feat(295), I1 =>  inp_feat(351), I2 =>  inp_feat(38), I3 =>  inp_feat(344), I4 =>  inp_feat(413), I5 =>  inp_feat(30), I6 =>  inp_feat(105), I7 =>  inp_feat(42)); 
C_24_S_3_L_7_inst : LUT8 generic map(INIT => "1111110100000101010000010000110111000001000101010011001101110100010010000000000000000000000000001000000000000000000000000000000011110000000100001111110101000101000000000001000100110011001101110010000000000000001000000000000000000000000100010000000000010001") port map( O =>C_24_S_3_L_7_out, I0 =>  inp_feat(98), I1 =>  inp_feat(506), I2 =>  inp_feat(445), I3 =>  inp_feat(242), I4 =>  inp_feat(40), I5 =>  inp_feat(51), I6 =>  inp_feat(300), I7 =>  inp_feat(322)); 
C_24_S_4_L_0_inst : LUT8 generic map(INIT => "0010100010101000101100001001000010101000100000001000000000000000001011100010101001000001101011111010001011101010101000001000101000001010000000000000000011000000100010101000000010000000100000000000000010000000000000001000000010000000100000001000000010000000") port map( O =>C_24_S_4_L_0_out, I0 =>  inp_feat(430), I1 =>  inp_feat(504), I2 =>  inp_feat(98), I3 =>  inp_feat(391), I4 =>  inp_feat(324), I5 =>  inp_feat(69), I6 =>  inp_feat(161), I7 =>  inp_feat(28)); 
C_24_S_4_L_1_inst : LUT8 generic map(INIT => "0010101011010010100110101110011110001110010000001010000011110000011000101100000000001100110000001111101111100000011101001011010011101110000000000000000000000000001110001110000011110000111000001010001000000000100011000100010011110010111100001111010010110100") port map( O =>C_24_S_4_L_1_out, I0 =>  inp_feat(41), I1 =>  inp_feat(82), I2 =>  inp_feat(506), I3 =>  inp_feat(328), I4 =>  inp_feat(161), I5 =>  inp_feat(114), I6 =>  inp_feat(413), I7 =>  inp_feat(83)); 
C_24_S_4_L_2_inst : LUT8 generic map(INIT => "0001000111101000000010100000100011011010001010001010001000100010000111111111010111111011111111011111111110111111101000101110111010101101110011001010100011001000101011001000001110011010001000101111100111111101111111111111111011011111111111110010111111111111") port map( O =>C_24_S_4_L_2_out, I0 =>  inp_feat(120), I1 =>  inp_feat(142), I2 =>  inp_feat(83), I3 =>  inp_feat(105), I4 =>  inp_feat(247), I5 =>  inp_feat(382), I6 =>  inp_feat(353), I7 =>  inp_feat(420)); 
C_24_S_4_L_3_inst : LUT8 generic map(INIT => "1111111010100000001110100010001010110010000000000011101000000010110110101010001001111010101010100010101000000000001110100000101011100000100000000010101000100010001010000000000000000000000000100001000000000000010110101010001000110000000000000010101000000010") port map( O =>C_24_S_4_L_3_out, I0 =>  inp_feat(309), I1 =>  inp_feat(295), I2 =>  inp_feat(344), I3 =>  inp_feat(30), I4 =>  inp_feat(296), I5 =>  inp_feat(238), I6 =>  inp_feat(478), I7 =>  inp_feat(303)); 
C_24_S_4_L_4_inst : LUT8 generic map(INIT => "1010101011101010111010001111111010000000001010001010101010101010100000101111101011101000111011110000001010001010000000001010000000101000101000000010010001100100000000000000000000000000000000000000000010000000001010000111000000000000000000000000000000000000") port map( O =>C_24_S_4_L_4_out, I0 =>  inp_feat(20), I1 =>  inp_feat(238), I2 =>  inp_feat(448), I3 =>  inp_feat(331), I4 =>  inp_feat(58), I5 =>  inp_feat(342), I6 =>  inp_feat(275), I7 =>  inp_feat(210)); 
C_24_S_4_L_5_inst : LUT8 generic map(INIT => "0110010101000000110000010000000010111011110011111100111000001110100000000000000010000000100000000000101000001000101000101010011001001000100011001000010000000000010000101000010011001110101011100000100000001000000000000000100000000000001000000010000000001010") port map( O =>C_24_S_4_L_5_out, I0 =>  inp_feat(365), I1 =>  inp_feat(327), I2 =>  inp_feat(180), I3 =>  inp_feat(99), I4 =>  inp_feat(74), I5 =>  inp_feat(351), I6 =>  inp_feat(417), I7 =>  inp_feat(31)); 
C_24_S_4_L_6_inst : LUT8 generic map(INIT => "0100101000101101111010101010111111001110110001001101000110101111100111010000110001000001100011000100111110001110100011111100111000000000000011000000000010001111000010100000001000001000100011010000000000000000000000000000000001001001000000001010110000001110") port map( O =>C_24_S_4_L_6_out, I0 =>  inp_feat(470), I1 =>  inp_feat(373), I2 =>  inp_feat(413), I3 =>  inp_feat(42), I4 =>  inp_feat(420), I5 =>  inp_feat(141), I6 =>  inp_feat(142), I7 =>  inp_feat(144)); 
C_24_S_4_L_7_inst : LUT8 generic map(INIT => "1111101011101010111111011111111110111010101000101111100000010001001000101010100101110010111100111111001010001000101111011111001100000000101101000000010111111101101000101110001000000000000010000001000001110001011001111111011000010010011110101111011111110111") port map( O =>C_24_S_4_L_7_out, I0 =>  inp_feat(120), I1 =>  inp_feat(362), I2 =>  inp_feat(500), I3 =>  inp_feat(316), I4 =>  inp_feat(477), I5 =>  inp_feat(382), I6 =>  inp_feat(29), I7 =>  inp_feat(52)); 
C_25_S_0_L_0_inst : LUT8 generic map(INIT => "0000000100000000001000000000001000000000000000000000000000000000000000000000100000100010100010100000000010000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000010000000100010101000101000000000000000000000000010001000") port map( O =>C_25_S_0_L_0_out, I0 =>  inp_feat(98), I1 =>  inp_feat(244), I2 =>  inp_feat(17), I3 =>  inp_feat(103), I4 =>  inp_feat(464), I5 =>  inp_feat(16), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_25_S_0_L_1_inst : LUT8 generic map(INIT => "1001000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_0_L_1_out, I0 =>  inp_feat(117), I1 =>  inp_feat(472), I2 =>  inp_feat(501), I3 =>  inp_feat(179), I4 =>  inp_feat(98), I5 =>  inp_feat(79), I6 =>  inp_feat(492), I7 =>  inp_feat(4)); 
C_25_S_0_L_2_inst : LUT8 generic map(INIT => "0000000011101000000000000000100000000000010010000000000000000000000000000000000000000000000000000000000010110000000000000000000010001000100010000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_0_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(92), I2 =>  inp_feat(29), I3 =>  inp_feat(249), I4 =>  inp_feat(479), I5 =>  inp_feat(218), I6 =>  inp_feat(293), I7 =>  inp_feat(229)); 
C_25_S_0_L_3_inst : LUT8 generic map(INIT => "0000000001110000000000000000000000000000000000000000000000000000100100001111000000010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_0_L_3_out, I0 =>  inp_feat(249), I1 =>  inp_feat(103), I2 =>  inp_feat(459), I3 =>  inp_feat(46), I4 =>  inp_feat(214), I5 =>  inp_feat(336), I6 =>  inp_feat(494), I7 =>  inp_feat(376)); 
C_25_S_0_L_4_inst : LUT8 generic map(INIT => "0000000011000000000000000000000001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000010000001100010000000000000000000000000000000000000000000000000001000000000000000000000000000000") port map( O =>C_25_S_0_L_4_out, I0 =>  inp_feat(75), I1 =>  inp_feat(336), I2 =>  inp_feat(239), I3 =>  inp_feat(29), I4 =>  inp_feat(158), I5 =>  inp_feat(340), I6 =>  inp_feat(332), I7 =>  inp_feat(117)); 
C_25_S_0_L_5_inst : LUT8 generic map(INIT => "0000100000000000000000000000000010001000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000010001000000000001000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_0_L_5_out, I0 =>  inp_feat(4), I1 =>  inp_feat(158), I2 =>  inp_feat(303), I3 =>  inp_feat(53), I4 =>  inp_feat(50), I5 =>  inp_feat(179), I6 =>  inp_feat(331), I7 =>  inp_feat(103)); 
C_25_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000110010000000000000000000000000000000000000000000110000000000000010000000010000000010000000000000010000000000000010000000000000001000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_25_S_0_L_6_out, I0 =>  inp_feat(195), I1 =>  inp_feat(263), I2 =>  inp_feat(493), I3 =>  inp_feat(381), I4 =>  inp_feat(157), I5 =>  inp_feat(50), I6 =>  inp_feat(249), I7 =>  inp_feat(159)); 
C_25_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000100000001000001010000000000000000000000000000000000000001000001010100010101000101000000000000010000000000010000000000010100000001000001010000000000000000000000000000000000000000000001010000000000000101000000000000000000000000000000000000000000000") port map( O =>C_25_S_0_L_7_out, I0 =>  inp_feat(462), I1 =>  inp_feat(460), I2 =>  inp_feat(445), I3 =>  inp_feat(117), I4 =>  inp_feat(157), I5 =>  inp_feat(50), I6 =>  inp_feat(249), I7 =>  inp_feat(144)); 
C_25_S_1_L_0_inst : LUT8 generic map(INIT => "0000000100000000001000000000001000000000000000000000000000000000000000000000100000100010100010100000000010000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000010000000100010101000101000000000000000000000000010001000") port map( O =>C_25_S_1_L_0_out, I0 =>  inp_feat(98), I1 =>  inp_feat(244), I2 =>  inp_feat(17), I3 =>  inp_feat(103), I4 =>  inp_feat(464), I5 =>  inp_feat(16), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_25_S_1_L_1_inst : LUT8 generic map(INIT => "1001000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_1_L_1_out, I0 =>  inp_feat(117), I1 =>  inp_feat(472), I2 =>  inp_feat(501), I3 =>  inp_feat(179), I4 =>  inp_feat(98), I5 =>  inp_feat(79), I6 =>  inp_feat(492), I7 =>  inp_feat(4)); 
C_25_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000101000000000100000000001100010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100011000000000000000000010011000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_1_L_2_out, I0 =>  inp_feat(15), I1 =>  inp_feat(200), I2 =>  inp_feat(464), I3 =>  inp_feat(71), I4 =>  inp_feat(36), I5 =>  inp_feat(29), I6 =>  inp_feat(336), I7 =>  inp_feat(256)); 
C_25_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000110000001000000000000000000000000000000000000000110100000100000011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_1_L_3_out, I0 =>  inp_feat(179), I1 =>  inp_feat(331), I2 =>  inp_feat(167), I3 =>  inp_feat(214), I4 =>  inp_feat(89), I5 =>  inp_feat(175), I6 =>  inp_feat(130), I7 =>  inp_feat(310)); 
C_25_S_1_L_4_inst : LUT8 generic map(INIT => "1000000010100000000000000000000010100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000110000000000000001000000000000001000000010000000000000000000000001000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_1_L_4_out, I0 =>  inp_feat(82), I1 =>  inp_feat(195), I2 =>  inp_feat(336), I3 =>  inp_feat(249), I4 =>  inp_feat(480), I5 =>  inp_feat(342), I6 =>  inp_feat(332), I7 =>  inp_feat(280)); 
C_25_S_1_L_5_inst : LUT8 generic map(INIT => "0001000101000000000100000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101011001000111010100000100000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_1_L_5_out, I0 =>  inp_feat(211), I1 =>  inp_feat(300), I2 =>  inp_feat(107), I3 =>  inp_feat(179), I4 =>  inp_feat(450), I5 =>  inp_feat(248), I6 =>  inp_feat(30), I7 =>  inp_feat(280)); 
C_25_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000001010000000000000110011000101100010100010000000000000000000000000000000000000000000000000000000000000000000000000000010001001100010110000000000000000100000000010101100000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_25_S_1_L_6_out, I0 =>  inp_feat(207), I1 =>  inp_feat(198), I2 =>  inp_feat(323), I3 =>  inp_feat(464), I4 =>  inp_feat(380), I5 =>  inp_feat(117), I6 =>  inp_feat(7), I7 =>  inp_feat(97)); 
C_25_S_1_L_7_inst : LUT8 generic map(INIT => "1110100000000000000010000000000010001000000010001000100000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_1_L_7_out, I0 =>  inp_feat(200), I1 =>  inp_feat(50), I2 =>  inp_feat(467), I3 =>  inp_feat(479), I4 =>  inp_feat(88), I5 =>  inp_feat(300), I6 =>  inp_feat(286), I7 =>  inp_feat(462)); 
C_25_S_2_L_0_inst : LUT8 generic map(INIT => "0000000100000000001000000000001000000000000000000000000000000000000000000000100000100010100010100000000010000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000010000000100010101000101000000000000000000000000010001000") port map( O =>C_25_S_2_L_0_out, I0 =>  inp_feat(98), I1 =>  inp_feat(244), I2 =>  inp_feat(17), I3 =>  inp_feat(103), I4 =>  inp_feat(464), I5 =>  inp_feat(16), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_25_S_2_L_1_inst : LUT8 generic map(INIT => "1001000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_2_L_1_out, I0 =>  inp_feat(117), I1 =>  inp_feat(472), I2 =>  inp_feat(501), I3 =>  inp_feat(179), I4 =>  inp_feat(98), I5 =>  inp_feat(79), I6 =>  inp_feat(492), I7 =>  inp_feat(4)); 
C_25_S_2_L_2_inst : LUT8 generic map(INIT => "0000010000000000011100000000000000000000000000000000000000000000001111000000000000110000000000000011000000000000000000000000000011001100000000000101000000000000000000000000000000000000000000001111110000000000001100000000000000101000000000000000000000000000") port map( O =>C_25_S_2_L_2_out, I0 =>  inp_feat(34), I1 =>  inp_feat(39), I2 =>  inp_feat(179), I3 =>  inp_feat(4), I4 =>  inp_feat(495), I5 =>  inp_feat(214), I6 =>  inp_feat(425), I7 =>  inp_feat(256)); 
C_25_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000110000000000000000000000000000000000000000000000110000100000000011000000010000000000000100000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_2_L_3_out, I0 =>  inp_feat(455), I1 =>  inp_feat(407), I2 =>  inp_feat(307), I3 =>  inp_feat(64), I4 =>  inp_feat(103), I5 =>  inp_feat(376), I6 =>  inp_feat(494), I7 =>  inp_feat(336)); 
C_25_S_2_L_4_inst : LUT8 generic map(INIT => "0010101000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001000010000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_2_L_4_out, I0 =>  inp_feat(286), I1 =>  inp_feat(250), I2 =>  inp_feat(95), I3 =>  inp_feat(354), I4 =>  inp_feat(204), I5 =>  inp_feat(117), I6 =>  inp_feat(30), I7 =>  inp_feat(464)); 
C_25_S_2_L_5_inst : LUT8 generic map(INIT => "0000100000001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100010001000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000") port map( O =>C_25_S_2_L_5_out, I0 =>  inp_feat(6), I1 =>  inp_feat(462), I2 =>  inp_feat(130), I3 =>  inp_feat(299), I4 =>  inp_feat(180), I5 =>  inp_feat(263), I6 =>  inp_feat(266), I7 =>  inp_feat(249)); 
C_25_S_2_L_6_inst : LUT8 generic map(INIT => "0010000000101000000000000000000010101010001000000000000000000000000000000000000000000000000000000010000000000000000000000000000010101010001010100000000000000000101010100010001000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_2_L_6_out, I0 =>  inp_feat(38), I1 =>  inp_feat(103), I2 =>  inp_feat(185), I3 =>  inp_feat(65), I4 =>  inp_feat(7), I5 =>  inp_feat(157), I6 =>  inp_feat(50), I7 =>  inp_feat(280)); 
C_25_S_2_L_7_inst : LUT8 generic map(INIT => "0010001100000010000000000000000010100010000000100000000000000000101010100000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000") port map( O =>C_25_S_2_L_7_out, I0 =>  inp_feat(53), I1 =>  inp_feat(464), I2 =>  inp_feat(249), I3 =>  inp_feat(270), I4 =>  inp_feat(92), I5 =>  inp_feat(259), I6 =>  inp_feat(280), I7 =>  inp_feat(332)); 
C_25_S_3_L_0_inst : LUT8 generic map(INIT => "0000000100000000001000000000001000000000000000000000000000000000000000000000100000100010100010100000000010000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000010000000100010101000101000000000000000000000000010001000") port map( O =>C_25_S_3_L_0_out, I0 =>  inp_feat(98), I1 =>  inp_feat(244), I2 =>  inp_feat(17), I3 =>  inp_feat(103), I4 =>  inp_feat(464), I5 =>  inp_feat(16), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_25_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000100000001000001010000000100000100000000000000010000000000000000010000000100000101000000000000000000000000000001000000000000000000000000000000000000000010000001000000000000000100000001000000000000000000000001000000010000000000000001000000010000000") port map( O =>C_25_S_3_L_1_out, I0 =>  inp_feat(472), I1 =>  inp_feat(144), I2 =>  inp_feat(474), I3 =>  inp_feat(249), I4 =>  inp_feat(464), I5 =>  inp_feat(117), I6 =>  inp_feat(157), I7 =>  inp_feat(452)); 
C_25_S_3_L_2_inst : LUT8 generic map(INIT => "0000000010010000000000001000000000000000101000010000000010000000101000001011000100000000000000000000000010100010000000000000000000100000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000100000000000000000000000") port map( O =>C_25_S_3_L_2_out, I0 =>  inp_feat(40), I1 =>  inp_feat(134), I2 =>  inp_feat(82), I3 =>  inp_feat(223), I4 =>  inp_feat(324), I5 =>  inp_feat(103), I6 =>  inp_feat(256), I7 =>  inp_feat(376)); 
C_25_S_3_L_3_inst : LUT8 generic map(INIT => "1000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_3_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(38), I2 =>  inp_feat(361), I3 =>  inp_feat(164), I4 =>  inp_feat(445), I5 =>  inp_feat(376), I6 =>  inp_feat(464), I7 =>  inp_feat(310)); 
C_25_S_3_L_4_inst : LUT8 generic map(INIT => "0000110000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_3_L_4_out, I0 =>  inp_feat(509), I1 =>  inp_feat(376), I2 =>  inp_feat(46), I3 =>  inp_feat(53), I4 =>  inp_feat(263), I5 =>  inp_feat(366), I6 =>  inp_feat(310), I7 =>  inp_feat(494)); 
C_25_S_3_L_5_inst : LUT8 generic map(INIT => "0001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000101000000000000000000000000000101010110000010000000000000000001000010100000000000000000000000010001000000000000000000000000000") port map( O =>C_25_S_3_L_5_out, I0 =>  inp_feat(71), I1 =>  inp_feat(207), I2 =>  inp_feat(179), I3 =>  inp_feat(98), I4 =>  inp_feat(176), I5 =>  inp_feat(274), I6 =>  inp_feat(485), I7 =>  inp_feat(509)); 
C_25_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000010000000000000000000000000000000000010000100000000000100000011100000000000000000000000000000000000000000010110000100000000001000000000000000000000000000000000000001100001011000010010000001100000000000000000000000000000000000000") port map( O =>C_25_S_3_L_6_out, I0 =>  inp_feat(95), I1 =>  inp_feat(179), I2 =>  inp_feat(117), I3 =>  inp_feat(280), I4 =>  inp_feat(437), I5 =>  inp_feat(442), I6 =>  inp_feat(509), I7 =>  inp_feat(249)); 
C_25_S_3_L_7_inst : LUT8 generic map(INIT => "0000100000111000010000000100000000000000000000000000000000000000010001011101010111001100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100010000000000000000000000000000000000000000000000") port map( O =>C_25_S_3_L_7_out, I0 =>  inp_feat(464), I1 =>  inp_feat(376), I2 =>  inp_feat(121), I3 =>  inp_feat(244), I4 =>  inp_feat(144), I5 =>  inp_feat(176), I6 =>  inp_feat(223), I7 =>  inp_feat(214)); 
C_25_S_4_L_0_inst : LUT8 generic map(INIT => "0000000100000000001000000000001000000000000000000000000000000000000000000000100000100010100010100000000010000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000010000000100010101000101000000000000000000000000010001000") port map( O =>C_25_S_4_L_0_out, I0 =>  inp_feat(98), I1 =>  inp_feat(244), I2 =>  inp_feat(17), I3 =>  inp_feat(103), I4 =>  inp_feat(464), I5 =>  inp_feat(16), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_25_S_4_L_1_inst : LUT8 generic map(INIT => "0000000100000011000101000000000000000000000000010000100000000001010100110001001100000000000000000001010100010011000100000000000100000000000100000000000000001001000000001000000000001000101000010000000100000000100100000100000000000000000000000001000000010000") port map( O =>C_25_S_4_L_1_out, I0 =>  inp_feat(249), I1 =>  inp_feat(464), I2 =>  inp_feat(228), I3 =>  inp_feat(244), I4 =>  inp_feat(117), I5 =>  inp_feat(399), I6 =>  inp_feat(18), I7 =>  inp_feat(452)); 
C_25_S_4_L_2_inst : LUT8 generic map(INIT => "1000110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_25_S_4_L_2_out, I0 =>  inp_feat(378), I1 =>  inp_feat(510), I2 =>  inp_feat(262), I3 =>  inp_feat(176), I4 =>  inp_feat(354), I5 =>  inp_feat(361), I6 =>  inp_feat(376), I7 =>  inp_feat(492)); 
C_25_S_4_L_3_inst : LUT8 generic map(INIT => "0000000001000000000000000100000011000000110000000000000001000000000000000000000000000000000000000100000010000000000000000000000001010000110000000000000011000000000000001100000000000000100000000000000000000000000000000000000000000000100000000000000000000000") port map( O =>C_25_S_4_L_3_out, I0 =>  inp_feat(509), I1 =>  inp_feat(307), I2 =>  inp_feat(200), I3 =>  inp_feat(178), I4 =>  inp_feat(214), I5 =>  inp_feat(103), I6 =>  inp_feat(376), I7 =>  inp_feat(256)); 
C_25_S_4_L_4_inst : LUT8 generic map(INIT => "0100110000000000000000000000001000001100000011000000000000000010000000000000000000000000000000000000000000000000000000000000000001001100000001001100110000001100010011000000110000000100000011100000000000000000000000000000000000000000000000000100010000000100") port map( O =>C_25_S_4_L_4_out, I0 =>  inp_feat(29), I1 =>  inp_feat(293), I2 =>  inp_feat(178), I3 =>  inp_feat(327), I4 =>  inp_feat(134), I5 =>  inp_feat(233), I6 =>  inp_feat(239), I7 =>  inp_feat(325)); 
C_25_S_4_L_5_inst : LUT8 generic map(INIT => "0111000001010000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000011000000000000000000000110000000100000001000000000000000000000000000000010000000000000000000000000000000000000000000000") port map( O =>C_25_S_4_L_5_out, I0 =>  inp_feat(244), I1 =>  inp_feat(93), I2 =>  inp_feat(474), I3 =>  inp_feat(376), I4 =>  inp_feat(53), I5 =>  inp_feat(450), I6 =>  inp_feat(378), I7 =>  inp_feat(179)); 
C_25_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000010100000000000000000000000000000001000000000100100000000000010110000000000001010000000000000101000000000000000000000000000000000000000000000100000000000001000000000000000100000000000000000101000000000000000100000000000001010001000000010") port map( O =>C_25_S_4_L_6_out, I0 =>  inp_feat(82), I1 =>  inp_feat(340), I2 =>  inp_feat(207), I3 =>  inp_feat(364), I4 =>  inp_feat(323), I5 =>  inp_feat(325), I6 =>  inp_feat(223), I7 =>  inp_feat(430)); 
C_25_S_4_L_7_inst : LUT8 generic map(INIT => "0000001000000111000000000000110000000000000000000000000000000000101000110000000000000000000000000000000000000000000000000000000011110111000001110000000000000000000000000000000000000000000000001011001100000000000000000000001000000000000000000000000000000000") port map( O =>C_25_S_4_L_7_out, I0 =>  inp_feat(305), I1 =>  inp_feat(52), I2 =>  inp_feat(134), I3 =>  inp_feat(14), I4 =>  inp_feat(53), I5 =>  inp_feat(310), I6 =>  inp_feat(77), I7 =>  inp_feat(299)); 
C_26_S_0_L_0_inst : LUT8 generic map(INIT => "1111110011100000101010001010000011111100111000001000100000000000101100001111000010100000101000000011000011000000000000000000000000000000000000000000100000000000101000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_0_L_0_out, I0 =>  inp_feat(25), I1 =>  inp_feat(479), I2 =>  inp_feat(464), I3 =>  inp_feat(69), I4 =>  inp_feat(161), I5 =>  inp_feat(390), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_26_S_0_L_1_inst : LUT8 generic map(INIT => "1101111111101010110001001100000011101111110010100001011111000000000011000000000000000100100000000000000000001010000100010100000000001100111010101100110011000000100000001110101000000000000000000000001000000000000000000000000000000000000000100000000000000000") port map( O =>C_26_S_0_L_1_out, I0 =>  inp_feat(331), I1 =>  inp_feat(29), I2 =>  inp_feat(407), I3 =>  inp_feat(479), I4 =>  inp_feat(438), I5 =>  inp_feat(139), I6 =>  inp_feat(300), I7 =>  inp_feat(211)); 
C_26_S_0_L_2_inst : LUT8 generic map(INIT => "1110100000100010110001000000100011001100100000001010110010000100110000000000000000000000000000001000000000000000000000000000000011101100001000101010110000000000111011000000000011101100100001001000000000000000000000000000000010000000000000001000000000000000") port map( O =>C_26_S_0_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(186), I2 =>  inp_feat(219), I3 =>  inp_feat(117), I4 =>  inp_feat(52), I5 =>  inp_feat(445), I6 =>  inp_feat(17), I7 =>  inp_feat(492)); 
C_26_S_0_L_3_inst : LUT8 generic map(INIT => "1111110011001100001010001000100010000000001000000000001000001000111110001111101000001000000010001011100010101010000000001000101000001001000010000000000000001000000000000000000000000000000000000101100000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_0_L_3_out, I0 =>  inp_feat(46), I1 =>  inp_feat(465), I2 =>  inp_feat(5), I3 =>  inp_feat(474), I4 =>  inp_feat(339), I5 =>  inp_feat(17), I6 =>  inp_feat(492), I7 =>  inp_feat(300)); 
C_26_S_0_L_4_inst : LUT8 generic map(INIT => "1011111100001000101011000010010010111000100000001000100000000000111111110000111111100100010001000000000000000000010000000000000000101000000000000000100000000000001000000000000000001000000000001000100000000000000000000000000000000000000000000000100000000000") port map( O =>C_26_S_0_L_4_out, I0 =>  inp_feat(509), I1 =>  inp_feat(183), I2 =>  inp_feat(176), I3 =>  inp_feat(300), I4 =>  inp_feat(98), I5 =>  inp_feat(113), I6 =>  inp_feat(493), I7 =>  inp_feat(223)); 
C_26_S_0_L_5_inst : LUT8 generic map(INIT => "0111100010100000100011111111110100001000000111001000100011101100111110001111000010001111111111110000000000000000000000000010110011000000000000001000100000000000000000000100000000001000000010001110000011100000100000000000000000000000000000000000000000001101") port map( O =>C_26_S_0_L_5_out, I0 =>  inp_feat(398), I1 =>  inp_feat(244), I2 =>  inp_feat(407), I3 =>  inp_feat(195), I4 =>  inp_feat(420), I5 =>  inp_feat(367), I6 =>  inp_feat(493), I7 =>  inp_feat(404)); 
C_26_S_0_L_6_inst : LUT8 generic map(INIT => "0010001010100010101100101010100010100000101000001111101110101000001000101010001000000010000000000000000000001000000000110000000010000000000000000011001100000000001000000000000000110011000000000001011100000000001100110000000000010001000000000011011100000000") port map( O =>C_26_S_0_L_6_out, I0 =>  inp_feat(464), I1 =>  inp_feat(331), I2 =>  inp_feat(274), I3 =>  inp_feat(358), I4 =>  inp_feat(376), I5 =>  inp_feat(298), I6 =>  inp_feat(17), I7 =>  inp_feat(341)); 
C_26_S_0_L_7_inst : LUT8 generic map(INIT => "0101111111111111111010001100110000001000010011000100110011011100111110001100010000001000010000001000000001000100000010000100010000000000110100000000000001000000000000000000000000000000110000001111000011010000000000000000000000000000000000000000000001000000") port map( O =>C_26_S_0_L_7_out, I0 =>  inp_feat(474), I1 =>  inp_feat(410), I2 =>  inp_feat(480), I3 =>  inp_feat(298), I4 =>  inp_feat(462), I5 =>  inp_feat(256), I6 =>  inp_feat(183), I7 =>  inp_feat(12)); 
C_26_S_1_L_0_inst : LUT8 generic map(INIT => "1111110011100000101010001010000011111100111000001000100000000000101100001111000010100000101000000011000011000000000000000000000000000000000000000000100000000000101000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_1_L_0_out, I0 =>  inp_feat(25), I1 =>  inp_feat(479), I2 =>  inp_feat(464), I3 =>  inp_feat(69), I4 =>  inp_feat(161), I5 =>  inp_feat(390), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_26_S_1_L_1_inst : LUT8 generic map(INIT => "1101111111101010110001001100000011101111110010100001011111000000000011000000000000000100100000000000000000001010000100010100000000001100111010101100110011000000100000001110101000000000000000000000001000000000000000000000000000000000000000100000000000000000") port map( O =>C_26_S_1_L_1_out, I0 =>  inp_feat(331), I1 =>  inp_feat(29), I2 =>  inp_feat(407), I3 =>  inp_feat(479), I4 =>  inp_feat(438), I5 =>  inp_feat(139), I6 =>  inp_feat(300), I7 =>  inp_feat(211)); 
C_26_S_1_L_2_inst : LUT8 generic map(INIT => "1111001011110000110000001001000010100010001000001100100001100000100000000111000000000000000000000010000000110000000000000000000010111010101100001100000011010000101010100011000011111000111100000000000001010000000000000000000000100000001100000011000001110000") port map( O =>C_26_S_1_L_2_out, I0 =>  inp_feat(222), I1 =>  inp_feat(125), I2 =>  inp_feat(18), I3 =>  inp_feat(302), I4 =>  inp_feat(52), I5 =>  inp_feat(445), I6 =>  inp_feat(17), I7 =>  inp_feat(492)); 
C_26_S_1_L_3_inst : LUT8 generic map(INIT => "1111001010110011000000000000000010101010101100001000101000000000100110001111100010001000100010000000000011110000000000000000000011001010110000000000000000000000100010101000000010000000100000001100000011000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_1_L_3_out, I0 =>  inp_feat(274), I1 =>  inp_feat(487), I2 =>  inp_feat(54), I3 =>  inp_feat(15), I4 =>  inp_feat(277), I5 =>  inp_feat(501), I6 =>  inp_feat(403), I7 =>  inp_feat(247)); 
C_26_S_1_L_4_inst : LUT8 generic map(INIT => "1111111100111010100000000000000011001100000000000000000000000000111111111101010100000000000000001100110000000000000000000000000011001100001000001100000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000") port map( O =>C_26_S_1_L_4_out, I0 =>  inp_feat(493), I1 =>  inp_feat(173), I2 =>  inp_feat(431), I3 =>  inp_feat(223), I4 =>  inp_feat(464), I5 =>  inp_feat(300), I6 =>  inp_feat(245), I7 =>  inp_feat(117)); 
C_26_S_1_L_5_inst : LUT8 generic map(INIT => "0110010000000000101010000000100011101100000010001010100000001000111011001010000010101000101010100001010000000000000000000000000010100000000000001010000000000000100000000000000010100000000000001010000000100000101000001010000000000000000000000000000000000000") port map( O =>C_26_S_1_L_5_out, I0 =>  inp_feat(63), I1 =>  inp_feat(69), I2 =>  inp_feat(381), I3 =>  inp_feat(277), I4 =>  inp_feat(480), I5 =>  inp_feat(403), I6 =>  inp_feat(501), I7 =>  inp_feat(318)); 
C_26_S_1_L_6_inst : LUT8 generic map(INIT => "0110111101001000111111010000000010101011000000001000100000000000111111110010001000010001000000001110111000100010000000000000000011101000001010000010000000100000000010000000000000000000000000000010000000110000001000000011000010000000000000000000000000000000") port map( O =>C_26_S_1_L_6_out, I0 =>  inp_feat(55), I1 =>  inp_feat(247), I2 =>  inp_feat(493), I3 =>  inp_feat(300), I4 =>  inp_feat(65), I5 =>  inp_feat(398), I6 =>  inp_feat(492), I7 =>  inp_feat(154)); 
C_26_S_1_L_7_inst : LUT8 generic map(INIT => "1011100010111010110111101110101001110000101000000111000010100010001010100110001000000010101010100000000000100000000000000000001010101010101000001000000011000000000000000000000011000000110000000010101000101010000000000000000000000000000000000000000000000000") port map( O =>C_26_S_1_L_7_out, I0 =>  inp_feat(117), I1 =>  inp_feat(239), I2 =>  inp_feat(322), I3 =>  inp_feat(307), I4 =>  inp_feat(381), I5 =>  inp_feat(93), I6 =>  inp_feat(274), I7 =>  inp_feat(260)); 
C_26_S_2_L_0_inst : LUT8 generic map(INIT => "1111110011100000101010001010000011111100111000001000100000000000101100001111000010100000101000000011000011000000000000000000000000000000000000000000100000000000101000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_2_L_0_out, I0 =>  inp_feat(25), I1 =>  inp_feat(479), I2 =>  inp_feat(464), I3 =>  inp_feat(69), I4 =>  inp_feat(161), I5 =>  inp_feat(390), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_26_S_2_L_1_inst : LUT8 generic map(INIT => "0001000011000000101100001000000011100000110100000000000011000000110100001000000010010000000100001110000010000000000000001000000011010000111111011011100011000000111000001100000010000000110000001001000000000000000100000000000010100000100000000000000000000000") port map( O =>C_26_S_2_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(54), I2 =>  inp_feat(299), I3 =>  inp_feat(442), I4 =>  inp_feat(501), I5 =>  inp_feat(264), I6 =>  inp_feat(79), I7 =>  inp_feat(272)); 
C_26_S_2_L_2_inst : LUT8 generic map(INIT => "1110111010111010100000001000101011001100111110100000000000001010000000001110001000000000000000101000000011101110000000000000000000011111101110101000001010001010000011000000100000001011000010100000001000000010000000001000101000000000000000000000000000000010") port map( O =>C_26_S_2_L_2_out, I0 =>  inp_feat(425), I1 =>  inp_feat(103), I2 =>  inp_feat(490), I3 =>  inp_feat(381), I4 =>  inp_feat(341), I5 =>  inp_feat(473), I6 =>  inp_feat(157), I7 =>  inp_feat(471)); 
C_26_S_2_L_3_inst : LUT8 generic map(INIT => "0111110100000101101011000000110011110000000000000010000010000000101011111000011110100010101010000010101000000000101000001010000011101100000000001010110010001100111110000000000010100000100000000010000000000000101000000000000000000000000000001010000010000000") port map( O =>C_26_S_2_L_3_out, I0 =>  inp_feat(502), I1 =>  inp_feat(408), I2 =>  inp_feat(438), I3 =>  inp_feat(97), I4 =>  inp_feat(435), I5 =>  inp_feat(493), I6 =>  inp_feat(336), I7 =>  inp_feat(57)); 
C_26_S_2_L_4_inst : LUT8 generic map(INIT => "1101010111110000110111000001000011010000111100000000000010111010111111011100000010001000101000100000000010100000101010001010001001000001010000000000000000000000000000000100000000000000000000000100000001000000000000001010000000000000000000000000000010101000") port map( O =>C_26_S_2_L_4_out, I0 =>  inp_feat(38), I1 =>  inp_feat(301), I2 =>  inp_feat(97), I3 =>  inp_feat(161), I4 =>  inp_feat(435), I5 =>  inp_feat(52), I6 =>  inp_feat(372), I7 =>  inp_feat(300)); 
C_26_S_2_L_5_inst : LUT8 generic map(INIT => "1010111000101010101011110001111100001000000000001001111100011001100011000000000010101110000000001100110000000000100011100000000000101010000000100000000000000000100000000000000000000000000000001010101000000000000000000000000010000000000000000000000000000000") port map( O =>C_26_S_2_L_5_out, I0 =>  inp_feat(464), I1 =>  inp_feat(438), I2 =>  inp_feat(331), I3 =>  inp_feat(25), I4 =>  inp_feat(347), I5 =>  inp_feat(52), I6 =>  inp_feat(161), I7 =>  inp_feat(267)); 
C_26_S_2_L_6_inst : LUT8 generic map(INIT => "1011110111001101110111001000100000001000000000001001100000000000110011000000100000001100100010001000100000000000100000000000000011110101000000000000110010001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000") port map( O =>C_26_S_2_L_6_out, I0 =>  inp_feat(435), I1 =>  inp_feat(509), I2 =>  inp_feat(331), I3 =>  inp_feat(235), I4 =>  inp_feat(378), I5 =>  inp_feat(256), I6 =>  inp_feat(47), I7 =>  inp_feat(404)); 
C_26_S_2_L_7_inst : LUT8 generic map(INIT => "1011101111110010001000001010001010111111111100110000000000101010100100001100000000000000000000001111111100110010000000000000000000000010101000000000000000000000100010000100000010000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_26_S_2_L_7_out, I0 =>  inp_feat(228), I1 =>  inp_feat(492), I2 =>  inp_feat(244), I3 =>  inp_feat(407), I4 =>  inp_feat(300), I5 =>  inp_feat(493), I6 =>  inp_feat(404), I7 =>  inp_feat(12)); 
C_26_S_3_L_0_inst : LUT8 generic map(INIT => "1111110011100000101010001010000011111100111000001000100000000000101100001111000010100000101000000011000011000000000000000000000000000000000000000000100000000000101000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_3_L_0_out, I0 =>  inp_feat(25), I1 =>  inp_feat(479), I2 =>  inp_feat(464), I3 =>  inp_feat(69), I4 =>  inp_feat(161), I5 =>  inp_feat(390), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_26_S_3_L_1_inst : LUT8 generic map(INIT => "0001000011000000101100001000000011100000110100000000000011000000110100001000000010010000000100001110000010000000000000001000000011010000111111011011100011000000111000001100000010000000110000001001000000000000000100000000000010100000100000000000000000000000") port map( O =>C_26_S_3_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(54), I2 =>  inp_feat(299), I3 =>  inp_feat(442), I4 =>  inp_feat(501), I5 =>  inp_feat(264), I6 =>  inp_feat(79), I7 =>  inp_feat(272)); 
C_26_S_3_L_2_inst : LUT8 generic map(INIT => "1111111111001000010010001000100011111000000010001000000010000000010101010000000000000000000000000000100000000000000000000000000001001101000010000100100010001000110010000000000010000000000000001101110100001000000000000000000000001000000000000000000000000000") port map( O =>C_26_S_3_L_2_out, I0 =>  inp_feat(183), I1 =>  inp_feat(25), I2 =>  inp_feat(492), I3 =>  inp_feat(179), I4 =>  inp_feat(342), I5 =>  inp_feat(117), I6 =>  inp_feat(341), I7 =>  inp_feat(471)); 
C_26_S_3_L_3_inst : LUT8 generic map(INIT => "1111110011010000100010001100000011110000000100001100000010000000111110101010000010101010000000000000000000000000000000000000000001100100001100000000000011100000010100001000000010000000000000001111011011110000101101101011000000000000000000000000000000000000") port map( O =>C_26_S_3_L_3_out, I0 =>  inp_feat(493), I1 =>  inp_feat(273), I2 =>  inp_feat(12), I3 =>  inp_feat(291), I4 =>  inp_feat(407), I5 =>  inp_feat(117), I6 =>  inp_feat(435), I7 =>  inp_feat(509)); 
C_26_S_3_L_4_inst : LUT8 generic map(INIT => "0111101101110000011110000000000011110000000000001111000001010000111100100000000010110000000000001111000000010000010100000100000001000000000010000000100000001000110000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_3_L_4_out, I0 =>  inp_feat(98), I1 =>  inp_feat(239), I2 =>  inp_feat(179), I3 =>  inp_feat(12), I4 =>  inp_feat(388), I5 =>  inp_feat(381), I6 =>  inp_feat(458), I7 =>  inp_feat(277)); 
C_26_S_3_L_5_inst : LUT8 generic map(INIT => "1111011001111011101000101010000011000010111000001010001000000000111000100000000011100000000000000000000000000000000000000000000011100000000000001000000000000000110000000100000000000000000000001010000000001010000000000000000000000000000000000000000000000000") port map( O =>C_26_S_3_L_5_out, I0 =>  inp_feat(339), I1 =>  inp_feat(364), I2 =>  inp_feat(156), I3 =>  inp_feat(99), I4 =>  inp_feat(141), I5 =>  inp_feat(277), I6 =>  inp_feat(458), I7 =>  inp_feat(117)); 
C_26_S_3_L_6_inst : LUT8 generic map(INIT => "0100110111111101111011001110111000000000110000001010100010001000111000001110100000100000001000000000000000000000001000000000000010111100110011001100110011001000101010000000000010001000000000001010000000000100000000000000000000000000000000000000000000000000") port map( O =>C_26_S_3_L_6_out, I0 =>  inp_feat(5), I1 =>  inp_feat(415), I2 =>  inp_feat(483), I3 =>  inp_feat(380), I4 =>  inp_feat(111), I5 =>  inp_feat(117), I6 =>  inp_feat(13), I7 =>  inp_feat(307)); 
C_26_S_3_L_7_inst : LUT8 generic map(INIT => "1111111011001010110010001000101000001000101010100000000000001010000001000000100010000000000000000000100010001010000010000000000011001100000000000000000000000000000000001000100000000000000000001110111010001000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_3_L_7_out, I0 =>  inp_feat(183), I1 =>  inp_feat(404), I2 =>  inp_feat(239), I3 =>  inp_feat(378), I4 =>  inp_feat(117), I5 =>  inp_feat(46), I6 =>  inp_feat(305), I7 =>  inp_feat(126)); 
C_26_S_4_L_0_inst : LUT8 generic map(INIT => "1111110011100000101010001010000011111100111000001000100000000000101100001111000010100000101000000011000011000000000000000000000000000000000000000000100000000000101000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_4_L_0_out, I0 =>  inp_feat(25), I1 =>  inp_feat(479), I2 =>  inp_feat(464), I3 =>  inp_feat(69), I4 =>  inp_feat(161), I5 =>  inp_feat(390), I6 =>  inp_feat(223), I7 =>  inp_feat(299)); 
C_26_S_4_L_1_inst : LUT8 generic map(INIT => "0001000011000000101100001000000011100000110100000000000011000000110100001000000010010000000100001110000010000000000000001000000011010000111111011011100011000000111000001100000010000000110000001001000000000000000100000000000010100000100000000000000000000000") port map( O =>C_26_S_4_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(54), I2 =>  inp_feat(299), I3 =>  inp_feat(442), I4 =>  inp_feat(501), I5 =>  inp_feat(264), I6 =>  inp_feat(79), I7 =>  inp_feat(272)); 
C_26_S_4_L_2_inst : LUT8 generic map(INIT => "1111110011001100110000001100010010001000000100000000100001100000110100000000000000000000000000001000100000000000000000000000000011100000100000001000000010000000100010000000000000000000010000001111000010000000000000000000000000001000000000000000000000000000") port map( O =>C_26_S_4_L_2_out, I0 =>  inp_feat(134), I1 =>  inp_feat(464), I2 =>  inp_feat(233), I3 =>  inp_feat(179), I4 =>  inp_feat(342), I5 =>  inp_feat(117), I6 =>  inp_feat(341), I7 =>  inp_feat(471)); 
C_26_S_4_L_3_inst : LUT8 generic map(INIT => "1000111010111011111100001111000000001100101100001011000010000000111111001010001010000000100000001010010010000000001000001000000011111010101010101010000000000000000000000000000000000000000000001111101010101010000000000000000000000000000000000000000000000000") port map( O =>C_26_S_4_L_3_out, I0 =>  inp_feat(145), I1 =>  inp_feat(494), I2 =>  inp_feat(152), I3 =>  inp_feat(158), I4 =>  inp_feat(502), I5 =>  inp_feat(117), I6 =>  inp_feat(493), I7 =>  inp_feat(435)); 
C_26_S_4_L_4_inst : LUT8 generic map(INIT => "1111101010001010000000000000000011111000011010100101000000000000111110000000101000000000000000101111100000100000111100000000000011110010000000100000000000100010101000001000000000110000000000001111101010001010101000101000101000100000000000000101000000000000") port map( O =>C_26_S_4_L_4_out, I0 =>  inp_feat(502), I1 =>  inp_feat(239), I2 =>  inp_feat(176), I3 =>  inp_feat(365), I4 =>  inp_feat(464), I5 =>  inp_feat(136), I6 =>  inp_feat(459), I7 =>  inp_feat(458)); 
C_26_S_4_L_5_inst : LUT8 generic map(INIT => "0100100000001000011111110000000011111010000000100000000000000010110010000000000011001100000000001100100000000000000000000000000011111101000001010111010100010101010111110000000101010111100101001100110001000000110001000000000000000000000000000000000000000000") port map( O =>C_26_S_4_L_5_out, I0 =>  inp_feat(98), I1 =>  inp_feat(381), I2 =>  inp_feat(474), I3 =>  inp_feat(12), I4 =>  inp_feat(201), I5 =>  inp_feat(455), I6 =>  inp_feat(318), I7 =>  inp_feat(307)); 
C_26_S_4_L_6_inst : LUT8 generic map(INIT => "1010110000001100111010000000000011001000100011001100000000000000101000100000000011001000000000000000000000000000000000000000000010100100100011001110100011000000100001001000000010100000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_26_S_4_L_6_out, I0 =>  inp_feat(97), I1 =>  inp_feat(93), I2 =>  inp_feat(455), I3 =>  inp_feat(256), I4 =>  inp_feat(420), I5 =>  inp_feat(47), I6 =>  inp_feat(404), I7 =>  inp_feat(480)); 
C_26_S_4_L_7_inst : LUT8 generic map(INIT => "0101011111100010111100111110000011000000111000001100000010000000100010101000000000100000101000001000000010000000110000000010000000001000100000001000000000000000000000000000000010100000101000000000000000000000101000001010000000000000000000001010000010100000") port map( O =>C_26_S_4_L_7_out, I0 =>  inp_feat(190), I1 =>  inp_feat(388), I2 =>  inp_feat(193), I3 =>  inp_feat(307), I4 =>  inp_feat(131), I5 =>  inp_feat(493), I6 =>  inp_feat(404), I7 =>  inp_feat(284)); 
C_27_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000100000000100000000000000010000000000000111000100000000001000000000000000000000000000000000000000000000101000000000000000000000000000001111000000000000000000000000000011110000000000000010000000000000") port map( O =>C_27_S_0_L_0_out, I0 =>  inp_feat(145), I1 =>  inp_feat(373), I2 =>  inp_feat(6), I3 =>  inp_feat(353), I4 =>  inp_feat(80), I5 =>  inp_feat(367), I6 =>  inp_feat(221), I7 =>  inp_feat(299)); 
C_27_S_0_L_1_inst : LUT8 generic map(INIT => "1110000110100000111100001000000001000000000000001101000000000000010111011000000011110010101000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_0_L_1_out, I0 =>  inp_feat(41), I1 =>  inp_feat(416), I2 =>  inp_feat(331), I3 =>  inp_feat(127), I4 =>  inp_feat(303), I5 =>  inp_feat(167), I6 =>  inp_feat(238), I7 =>  inp_feat(405)); 
C_27_S_0_L_2_inst : LUT8 generic map(INIT => "1101001000000000000000000000000001100000000000000000000000000000111100101000000010000000000000001111000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_27_S_0_L_2_out, I0 =>  inp_feat(179), I1 =>  inp_feat(436), I2 =>  inp_feat(508), I3 =>  inp_feat(100), I4 =>  inp_feat(251), I5 =>  inp_feat(413), I6 =>  inp_feat(29), I7 =>  inp_feat(148)); 
C_27_S_0_L_3_inst : LUT8 generic map(INIT => "0110011011111010000010000100100010100000000110000000000000000000000000001000000000000000000000000000000000000000000000000000000010100000110100000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_0_L_3_out, I0 =>  inp_feat(478), I1 =>  inp_feat(291), I2 =>  inp_feat(259), I3 =>  inp_feat(29), I4 =>  inp_feat(362), I5 =>  inp_feat(290), I6 =>  inp_feat(83), I7 =>  inp_feat(328)); 
C_27_S_0_L_4_inst : LUT8 generic map(INIT => "0100000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000011110100000000000001111100000000111100000000000000000000000000000100000001000000000000001000000000000000010000000000000000000000") port map( O =>C_27_S_0_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(283), I2 =>  inp_feat(105), I3 =>  inp_feat(324), I4 =>  inp_feat(310), I5 =>  inp_feat(276), I6 =>  inp_feat(506), I7 =>  inp_feat(509)); 
C_27_S_0_L_5_inst : LUT8 generic map(INIT => "1000101010000000000000000000000000000011100000000000000000000000101011110010000000000000001000000000000000000000000000000000000000110001100000000010001000000000000100001000000000100000000000000000000000100000000000000000000000000010000000000000001100100000") port map( O =>C_27_S_0_L_5_out, I0 =>  inp_feat(7), I1 =>  inp_feat(218), I2 =>  inp_feat(302), I3 =>  inp_feat(317), I4 =>  inp_feat(492), I5 =>  inp_feat(493), I6 =>  inp_feat(134), I7 =>  inp_feat(247)); 
C_27_S_0_L_6_inst : LUT8 generic map(INIT => "0100000010000000010000011101000000000000010000000100000001000101000000000000000000000000000001000000000001000000000001000000000010000000110000001100000011000000010001000000000000000000000000000100110001000100000000000000000001000000000000000000000000000100") port map( O =>C_27_S_0_L_6_out, I0 =>  inp_feat(509), I1 =>  inp_feat(444), I2 =>  inp_feat(98), I3 =>  inp_feat(97), I4 =>  inp_feat(24), I5 =>  inp_feat(473), I6 =>  inp_feat(60), I7 =>  inp_feat(460)); 
C_27_S_0_L_7_inst : LUT8 generic map(INIT => "1111001000100000100100100010000011100000101000000100000000000000000000000000000000100000000000000000000000001010000000000000000011100000001100000010000010110000101000001010000000000000101100000000000000110000000000000000000000001000000000100000001000000100") port map( O =>C_27_S_0_L_7_out, I0 =>  inp_feat(420), I1 =>  inp_feat(373), I2 =>  inp_feat(477), I3 =>  inp_feat(470), I4 =>  inp_feat(362), I5 =>  inp_feat(116), I6 =>  inp_feat(148), I7 =>  inp_feat(144)); 
C_27_S_1_L_0_inst : LUT8 generic map(INIT => "0010100000100000000000000000000010100000010000000001100100010000000000000000000000000000000000000000000000000000000000000000000010101110110000000000000000000000111100010000000000000000000000000000001100000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_1_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(301), I2 =>  inp_feat(141), I3 =>  inp_feat(328), I4 =>  inp_feat(105), I5 =>  inp_feat(303), I6 =>  inp_feat(405), I7 =>  inp_feat(210)); 
C_27_S_1_L_1_inst : LUT8 generic map(INIT => "1000000001000000100000000000000000000000000000000010000010010000000000000000010000000000000000000000000000000000000000000000000011000000110011001000000000000000000001000000000000000000000000000000001010000100000000000000000010000000000000000000000000000000") port map( O =>C_27_S_1_L_1_out, I0 =>  inp_feat(109), I1 =>  inp_feat(413), I2 =>  inp_feat(475), I3 =>  inp_feat(449), I4 =>  inp_feat(34), I5 =>  inp_feat(324), I6 =>  inp_feat(158), I7 =>  inp_feat(340)); 
C_27_S_1_L_2_inst : LUT8 generic map(INIT => "1010000000000000001100000010000000100000000011000010000000000000000000000000000000010000000000000001000000000000110100000000000000100000000000001010100000000000000000000000100011111000000000000000000000000000000000000000000000000000000000000100100000000000") port map( O =>C_27_S_1_L_2_out, I0 =>  inp_feat(451), I1 =>  inp_feat(464), I2 =>  inp_feat(224), I3 =>  inp_feat(195), I4 =>  inp_feat(178), I5 =>  inp_feat(373), I6 =>  inp_feat(331), I7 =>  inp_feat(95)); 
C_27_S_1_L_3_inst : LUT8 generic map(INIT => "0010000000010000111000000011000001000010011100001010000011110000101000000000000010010010001010000000000001010000101000001000001000000000000000000110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_1_L_3_out, I0 =>  inp_feat(451), I1 =>  inp_feat(221), I2 =>  inp_feat(83), I3 =>  inp_feat(380), I4 =>  inp_feat(52), I5 =>  inp_feat(30), I6 =>  inp_feat(141), I7 =>  inp_feat(506)); 
C_27_S_1_L_4_inst : LUT8 generic map(INIT => "1110111111011100011110000000000001010100010100110000100000000000110000001100000000000000000000001100000011110000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000010011000000000000000000010000000011000000100000000000000") port map( O =>C_27_S_1_L_4_out, I0 =>  inp_feat(373), I1 =>  inp_feat(362), I2 =>  inp_feat(316), I3 =>  inp_feat(144), I4 =>  inp_feat(413), I5 =>  inp_feat(470), I6 =>  inp_feat(116), I7 =>  inp_feat(148)); 
C_27_S_1_L_5_inst : LUT8 generic map(INIT => "0000010011101000011000000100000001000000110000001100011011000000000000000000000000000000000000000000000000000000000000000000000001110011011100001100001000000000000001001011110000000000010000000000000001100000000000000000000001000000110010000001000000000000") port map( O =>C_27_S_1_L_5_out, I0 =>  inp_feat(373), I1 =>  inp_feat(82), I2 =>  inp_feat(420), I3 =>  inp_feat(144), I4 =>  inp_feat(303), I5 =>  inp_feat(470), I6 =>  inp_feat(353), I7 =>  inp_feat(449)); 
C_27_S_1_L_6_inst : LUT8 generic map(INIT => "0100000011111100000000100011000100100000010111000000000000000100000000000000010000000000000000001000000000010101000000000000000011110000111100001100000011000000110100000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_1_L_6_out, I0 =>  inp_feat(41), I1 =>  inp_feat(58), I2 =>  inp_feat(161), I3 =>  inp_feat(52), I4 =>  inp_feat(416), I5 =>  inp_feat(247), I6 =>  inp_feat(273), I7 =>  inp_feat(18)); 
C_27_S_1_L_7_inst : LUT8 generic map(INIT => "1001000000000000000000000000110000000000000000001010000010000000011110100000100011001001100000000000000000000000000000010000000010000000000000000001000010011000000000000000000010000000100000000000000000000000100000001000000000000000000000000000000010001100") port map( O =>C_27_S_1_L_7_out, I0 =>  inp_feat(480), I1 =>  inp_feat(290), I2 =>  inp_feat(74), I3 =>  inp_feat(362), I4 =>  inp_feat(142), I5 =>  inp_feat(153), I6 =>  inp_feat(31), I7 =>  inp_feat(339)); 
C_27_S_2_L_0_inst : LUT8 generic map(INIT => "0000000100000000000010100000110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010100010110010101010010000001010100010001100100010001000000000100000000000001100110000000000001001000010011010000000100000") port map( O =>C_27_S_2_L_0_out, I0 =>  inp_feat(74), I1 =>  inp_feat(221), I2 =>  inp_feat(509), I3 =>  inp_feat(420), I4 =>  inp_feat(339), I5 =>  inp_feat(470), I6 =>  inp_feat(182), I7 =>  inp_feat(29)); 
C_27_S_2_L_1_inst : LUT8 generic map(INIT => "1101110000000100111110001000010011001110000001001001000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_2_L_1_out, I0 =>  inp_feat(308), I1 =>  inp_feat(247), I2 =>  inp_feat(18), I3 =>  inp_feat(183), I4 =>  inp_feat(478), I5 =>  inp_feat(491), I6 =>  inp_feat(508), I7 =>  inp_feat(331)); 
C_27_S_2_L_2_inst : LUT8 generic map(INIT => "0000100010111000010010001000101000000000000010000000010000000000100010000000100010001100100011010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000") port map( O =>C_27_S_2_L_2_out, I0 =>  inp_feat(161), I1 =>  inp_feat(273), I2 =>  inp_feat(509), I3 =>  inp_feat(15), I4 =>  inp_feat(29), I5 =>  inp_feat(309), I6 =>  inp_feat(130), I7 =>  inp_feat(100)); 
C_27_S_2_L_3_inst : LUT8 generic map(INIT => "0000001000000001101010011010000000000000000000000000000000000000000000000000001000110000111010000000000010000000100000001000100010010011101100001010001010100000000000000000000000000000000000000001100000001000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_2_L_3_out, I0 =>  inp_feat(380), I1 =>  inp_feat(228), I2 =>  inp_feat(4), I3 =>  inp_feat(256), I4 =>  inp_feat(130), I5 =>  inp_feat(100), I6 =>  inp_feat(224), I7 =>  inp_feat(178)); 
C_27_S_2_L_4_inst : LUT8 generic map(INIT => "1000110100000000001000000100000010000101001000000100000000000000000101000000000000000000000000001010100000000000000001000000000011110100000000000001001000000000000000000000000000000000010000000011001000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_2_L_4_out, I0 =>  inp_feat(41), I1 =>  inp_feat(90), I2 =>  inp_feat(504), I3 =>  inp_feat(86), I4 =>  inp_feat(449), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(238)); 
C_27_S_2_L_5_inst : LUT8 generic map(INIT => "1100000001000000010011000000000000000100000000000100010000000000000000000000000000000000010001000100000000000000000000000100000011000100000000001100110101000100000000000000000001001000000000000000000001000001010001000100000000000000010000001100010000000100") port map( O =>C_27_S_2_L_5_out, I0 =>  inp_feat(29), I1 =>  inp_feat(6), I2 =>  inp_feat(382), I3 =>  inp_feat(62), I4 =>  inp_feat(308), I5 =>  inp_feat(316), I6 =>  inp_feat(385), I7 =>  inp_feat(373)); 
C_27_S_2_L_6_inst : LUT8 generic map(INIT => "1011011100001111111010100001000000000000000000000000000000000000010010001000111010011000000000100000000000000000000000000000000000001000000010000000000000000000000000000000000000000000101000000000000110001110000000001011100000000000000000000000000010000000") port map( O =>C_27_S_2_L_6_out, I0 =>  inp_feat(316), I1 =>  inp_feat(420), I2 =>  inp_feat(467), I3 =>  inp_feat(38), I4 =>  inp_feat(95), I5 =>  inp_feat(148), I6 =>  inp_feat(259), I7 =>  inp_feat(354)); 
C_27_S_2_L_7_inst : LUT8 generic map(INIT => "0010111100000000010001000000100010001100000000101100000000000000100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_2_L_7_out, I0 =>  inp_feat(344), I1 =>  inp_feat(127), I2 =>  inp_feat(238), I3 =>  inp_feat(477), I4 =>  inp_feat(364), I5 =>  inp_feat(37), I6 =>  inp_feat(410), I7 =>  inp_feat(69)); 
C_27_S_3_L_0_inst : LUT8 generic map(INIT => "1010100000000001000000000010100010010000111000000000000010000000000000000010000000000000000000001010000000100000000000000000000000000000001000000000000010000000100000000010110000000000110010000010000000000000000000000000000010100010101001000000000010000100") port map( O =>C_27_S_3_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(178), I2 =>  inp_feat(422), I3 =>  inp_feat(41), I4 =>  inp_feat(493), I5 =>  inp_feat(29), I6 =>  inp_feat(233), I7 =>  inp_feat(346)); 
C_27_S_3_L_1_inst : LUT8 generic map(INIT => "1100110001010000100000000000000000000000000000000010000000000000111011100000000010001000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000001010110000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_3_L_1_out, I0 =>  inp_feat(365), I1 =>  inp_feat(351), I2 =>  inp_feat(350), I3 =>  inp_feat(286), I4 =>  inp_feat(125), I5 =>  inp_feat(69), I6 =>  inp_feat(18), I7 =>  inp_feat(480)); 
C_27_S_3_L_2_inst : LUT8 generic map(INIT => "0000001000101000101000001010110001101000001000111010000010101000111000011011011011100000101000000000000000111011100000001010001100000000000010000000000000000000000000000000000010100000000000000000000000000000000000001000000000000000000000000010010000000000") port map( O =>C_27_S_3_L_2_out, I0 =>  inp_feat(420), I1 =>  inp_feat(373), I2 =>  inp_feat(362), I3 =>  inp_feat(259), I4 =>  inp_feat(116), I5 =>  inp_feat(470), I6 =>  inp_feat(120), I7 =>  inp_feat(353)); 
C_27_S_3_L_3_inst : LUT8 generic map(INIT => "1011000000001000000000000000000010101000000000000000100000000000001000000000000000000000000000001011001000001010000000000000000000000010101000000001000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_3_L_3_out, I0 =>  inp_feat(6), I1 =>  inp_feat(373), I2 =>  inp_feat(316), I3 =>  inp_feat(111), I4 =>  inp_feat(477), I5 =>  inp_feat(238), I6 =>  inp_feat(331), I7 =>  inp_feat(62)); 
C_27_S_3_L_4_inst : LUT8 generic map(INIT => "1100100000101000001110000000000000001000001000000000100000000000000000001000000010101110000010000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000") port map( O =>C_27_S_3_L_4_out, I0 =>  inp_feat(57), I1 =>  inp_feat(3), I2 =>  inp_feat(291), I3 =>  inp_feat(115), I4 =>  inp_feat(399), I5 =>  inp_feat(506), I6 =>  inp_feat(256), I7 =>  inp_feat(403)); 
C_27_S_3_L_5_inst : LUT8 generic map(INIT => "0110111000001110001000100000010011101010000000000000110000000000000000000000000000000000000000000100100000000000000000000000000000001000001000000000000000000100000001000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000") port map( O =>C_27_S_3_L_5_out, I0 =>  inp_feat(478), I1 =>  inp_feat(277), I2 =>  inp_feat(303), I3 =>  inp_feat(66), I4 =>  inp_feat(479), I5 =>  inp_feat(151), I6 =>  inp_feat(309), I7 =>  inp_feat(87)); 
C_27_S_3_L_6_inst : LUT8 generic map(INIT => "0000111000010000000000000000000000100100000010000100000000000000000000000000000000000000000000000010010000001000100000000000000010001110101010100110000010100000111000001000000000000000001000000000001000000010000000000000100000000000100000001000001000000000") port map( O =>C_27_S_3_L_6_out, I0 =>  inp_feat(493), I1 =>  inp_feat(238), I2 =>  inp_feat(74), I3 =>  inp_feat(449), I4 =>  inp_feat(382), I5 =>  inp_feat(303), I6 =>  inp_feat(413), I7 =>  inp_feat(228)); 
C_27_S_3_L_7_inst : LUT8 generic map(INIT => "1000010010000001010001100000010001000100000001001010110001000000010001000000000001000100000000000100010000000000110001100010000000000000000001000000000000000000101000000000000010000001000000001000000000000000000010100000100011000000000000000000000000100000") port map( O =>C_27_S_3_L_7_out, I0 =>  inp_feat(221), I1 =>  inp_feat(344), I2 =>  inp_feat(340), I3 =>  inp_feat(504), I4 =>  inp_feat(177), I5 =>  inp_feat(238), I6 =>  inp_feat(275), I7 =>  inp_feat(290)); 
C_27_S_4_L_0_inst : LUT8 generic map(INIT => "1010100010101000101000000000100000000000000010000000000000000000100000001000101010100010100000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_27_S_4_L_0_out, I0 =>  inp_feat(508), I1 =>  inp_feat(50), I2 =>  inp_feat(351), I3 =>  inp_feat(277), I4 =>  inp_feat(478), I5 =>  inp_feat(477), I6 =>  inp_feat(320), I7 =>  inp_feat(161)); 
C_27_S_4_L_1_inst : LUT8 generic map(INIT => "1000011000001100000001000000000010110000010111000000000000000000000001000000011000000010000000000000000001101100000000000000000011001100100010001000000010001000100000001000000000000000000000000000000011001100000000000000000000000000010000000000000000000000") port map( O =>C_27_S_4_L_1_out, I0 =>  inp_feat(238), I1 =>  inp_feat(74), I2 =>  inp_feat(373), I3 =>  inp_feat(162), I4 =>  inp_feat(477), I5 =>  inp_feat(475), I6 =>  inp_feat(362), I7 =>  inp_feat(116)); 
C_27_S_4_L_2_inst : LUT8 generic map(INIT => "0111110001010000001010010000001000000000000000000000001010000000101000001111000000110000000100000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000100010000010110000000000110000000000000000000010001010101010001010") port map( O =>C_27_S_4_L_2_out, I0 =>  inp_feat(413), I1 =>  inp_feat(221), I2 =>  inp_feat(449), I3 =>  inp_feat(420), I4 =>  inp_feat(106), I5 =>  inp_feat(331), I6 =>  inp_feat(509), I7 =>  inp_feat(451)); 
C_27_S_4_L_3_inst : LUT8 generic map(INIT => "0011100011010000001111011000000000000000000000000001000100100000101100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000") port map( O =>C_27_S_4_L_3_out, I0 =>  inp_feat(97), I1 =>  inp_feat(242), I2 =>  inp_feat(216), I3 =>  inp_feat(177), I4 =>  inp_feat(478), I5 =>  inp_feat(7), I6 =>  inp_feat(238), I7 =>  inp_feat(482)); 
C_27_S_4_L_4_inst : LUT8 generic map(INIT => "0100100000001010100000000000000001000000101000000000000000000000110010000000000000000000000000000000100000000000000000000000110000101000000000000000000000000000011000100000001000000000000000001000101000001000100000000000000000100010000000100000000000000110") port map( O =>C_27_S_4_L_4_out, I0 =>  inp_feat(504), I1 =>  inp_feat(86), I2 =>  inp_feat(387), I3 =>  inp_feat(5), I4 =>  inp_feat(87), I5 =>  inp_feat(376), I6 =>  inp_feat(256), I7 =>  inp_feat(43)); 
C_27_S_4_L_5_inst : LUT8 generic map(INIT => "0000001010100001000000101010001000111010000010010000000000000000000000001000011000000000000000100100001000110011001100000001000000100000011000000000000010100010010001011110000100000000101000000100000010110101000000001010000000000001101001110000000010100000") port map( O =>C_27_S_4_L_5_out, I0 =>  inp_feat(141), I1 =>  inp_feat(52), I2 =>  inp_feat(420), I3 =>  inp_feat(221), I4 =>  inp_feat(294), I5 =>  inp_feat(308), I6 =>  inp_feat(470), I7 =>  inp_feat(95)); 
C_27_S_4_L_6_inst : LUT8 generic map(INIT => "0100101000000000110001000100000011010010000000000100000000000000000000000000000000000000000100001000000100000000000000010000000000000100000000000000000001010000000001000000010000000000000000000011000000010000001000000000001000100000000000000000000000000000") port map( O =>C_27_S_4_L_6_out, I0 =>  inp_feat(365), I1 =>  inp_feat(413), I2 =>  inp_feat(504), I3 =>  inp_feat(344), I4 =>  inp_feat(177), I5 =>  inp_feat(478), I6 =>  inp_feat(87), I7 =>  inp_feat(316)); 
C_27_S_4_L_7_inst : LUT8 generic map(INIT => "1110011010001110000000001001000100010010000000000111010000100000110000000000000000000000000000000000000000000000000000000000000010000000000000001010000000000000000000000000000000000000000000001010000000000000001000000000000000000000000000001010000000000000") port map( O =>C_27_S_4_L_7_out, I0 =>  inp_feat(398), I1 =>  inp_feat(244), I2 =>  inp_feat(296), I3 =>  inp_feat(205), I4 =>  inp_feat(262), I5 =>  inp_feat(445), I6 =>  inp_feat(74), I7 =>  inp_feat(14)); 
C_28_S_0_L_0_inst : LUT8 generic map(INIT => "0100000000000000000000000000000000000100000000000000000000000000011111110000000000000000000000000000110000000000000000000000000000001111000000000000001000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_0_L_0_out, I0 =>  inp_feat(256), I1 =>  inp_feat(180), I2 =>  inp_feat(494), I3 =>  inp_feat(98), I4 =>  inp_feat(331), I5 =>  inp_feat(372), I6 =>  inp_feat(157), I7 =>  inp_feat(299)); 
C_28_S_0_L_1_inst : LUT8 generic map(INIT => "1110101110010001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101100100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_0_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(18), I2 =>  inp_feat(295), I3 =>  inp_feat(504), I4 =>  inp_feat(361), I5 =>  inp_feat(403), I6 =>  inp_feat(405), I7 =>  inp_feat(210)); 
C_28_S_0_L_2_inst : LUT8 generic map(INIT => "0010001111111100000000001000000011100000111100000000000000000000000000000000000000000000100000000101000000000000000000000000000011100000111100000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_0_L_2_out, I0 =>  inp_feat(323), I1 =>  inp_feat(52), I2 =>  inp_feat(378), I3 =>  inp_feat(223), I4 =>  inp_feat(167), I5 =>  inp_feat(238), I6 =>  inp_feat(413), I7 =>  inp_feat(144)); 
C_28_S_0_L_3_inst : LUT8 generic map(INIT => "0111111100000000000001000000000010000000000000010000000000000000010000010000000000000001000000000000000000000000000000000000000011110111000000000000000000000000000100010000000100000000000000000000001010000000000000100000000000000001000000000000000000000000") port map( O =>C_28_S_0_L_3_out, I0 =>  inp_feat(394), I1 =>  inp_feat(29), I2 =>  inp_feat(509), I3 =>  inp_feat(331), I4 =>  inp_feat(478), I5 =>  inp_feat(283), I6 =>  inp_feat(420), I7 =>  inp_feat(373)); 
C_28_S_0_L_4_inst : LUT8 generic map(INIT => "1110010010000000001000000000000000000001000000000000000000000000110000001000000000001000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000001001000100000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_0_L_4_out, I0 =>  inp_feat(346), I1 =>  inp_feat(86), I2 =>  inp_feat(435), I3 =>  inp_feat(295), I4 =>  inp_feat(344), I5 =>  inp_feat(506), I6 =>  inp_feat(256), I7 =>  inp_feat(247)); 
C_28_S_0_L_5_inst : LUT8 generic map(INIT => "1000100010000000100001001101000110000000000000001000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100") port map( O =>C_28_S_0_L_5_out, I0 =>  inp_feat(141), I1 =>  inp_feat(331), I2 =>  inp_feat(413), I3 =>  inp_feat(177), I4 =>  inp_feat(420), I5 =>  inp_feat(342), I6 =>  inp_feat(80), I7 =>  inp_feat(290)); 
C_28_S_0_L_6_inst : LUT8 generic map(INIT => "1000100000000001000000001000100000100000000000000000000000000000101000101000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001011000000000000001000000011000000000000000000000000000000000000") port map( O =>C_28_S_0_L_6_out, I0 =>  inp_feat(98), I1 =>  inp_feat(420), I2 =>  inp_feat(344), I3 =>  inp_feat(413), I4 =>  inp_feat(408), I5 =>  inp_feat(506), I6 =>  inp_feat(256), I7 =>  inp_feat(247)); 
C_28_S_0_L_7_inst : LUT8 generic map(INIT => "0000101000001000000010000000100000000000000000000000000000000000100010000000000000000000100000001011000000000000000000000000000011001000000000001000110000001010000000000000000000000000000000001100100000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_0_L_7_out, I0 =>  inp_feat(331), I1 =>  inp_feat(23), I2 =>  inp_feat(97), I3 =>  inp_feat(273), I4 =>  inp_feat(478), I5 =>  inp_feat(287), I6 =>  inp_feat(54), I7 =>  inp_feat(367)); 
C_28_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000110000000000000001000000000000001100000000000000000000000000000000100100010000000000000000000000100000000000000011001010100000001100000000000000100010000000000011000000000000000000000000000000000000000000000000001000100010000000000000000000") port map( O =>C_28_S_1_L_0_out, I0 =>  inp_feat(471), I1 =>  inp_feat(344), I2 =>  inp_feat(331), I3 =>  inp_feat(347), I4 =>  inp_feat(25), I5 =>  inp_feat(275), I6 =>  inp_feat(420), I7 =>  inp_feat(335)); 
C_28_S_1_L_1_inst : LUT8 generic map(INIT => "0000110101001000010001110100000000000111000000000000000000000000000000000000000000010010000000000000000000000000000000000000000011000100000000000100010100000100000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000") port map( O =>C_28_S_1_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(478), I2 =>  inp_feat(356), I3 =>  inp_feat(281), I4 =>  inp_feat(256), I5 =>  inp_feat(506), I6 =>  inp_feat(232), I7 =>  inp_feat(460)); 
C_28_S_1_L_2_inst : LUT8 generic map(INIT => "1100101000000000100010001000000010001000000000001000100010000000000000000000000000001000000010001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_1_L_2_out, I0 =>  inp_feat(152), I1 =>  inp_feat(98), I2 =>  inp_feat(484), I3 =>  inp_feat(447), I4 =>  inp_feat(18), I5 =>  inp_feat(346), I6 =>  inp_feat(217), I7 =>  inp_feat(474)); 
C_28_S_1_L_3_inst : LUT8 generic map(INIT => "1010010001100100100000000000000011100000010000000010000000000000100000000000000000000000000000001100000100100101000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000100000000000000000000000001000100000000100000001000000") port map( O =>C_28_S_1_L_3_out, I0 =>  inp_feat(380), I1 =>  inp_feat(420), I2 =>  inp_feat(83), I3 =>  inp_feat(362), I4 =>  inp_feat(413), I5 =>  inp_feat(373), I6 =>  inp_feat(42), I7 =>  inp_feat(477)); 
C_28_S_1_L_4_inst : LUT8 generic map(INIT => "0000101010100010011011100010001000000000010010001111101110000100001000101000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_1_L_4_out, I0 =>  inp_feat(161), I1 =>  inp_feat(116), I2 =>  inp_feat(120), I3 =>  inp_feat(145), I4 =>  inp_feat(259), I5 =>  inp_feat(362), I6 =>  inp_feat(477), I7 =>  inp_feat(474)); 
C_28_S_1_L_5_inst : LUT8 generic map(INIT => "0000110000000000010011000000000000111100000000001100010001000000000001001000000011001111000011000100010000000000010001000000000000000000000000000000010000000000000000000000000000000000000000000000110100000000010000100000010000000000000000000000000000000000") port map( O =>C_28_S_1_L_5_out, I0 =>  inp_feat(221), I1 =>  inp_feat(290), I2 =>  inp_feat(367), I3 =>  inp_feat(82), I4 =>  inp_feat(41), I5 =>  inp_feat(277), I6 =>  inp_feat(19), I7 =>  inp_feat(62)); 
C_28_S_1_L_6_inst : LUT8 generic map(INIT => "0100000000100000110010000000101000001000000000000000000000000000000000000000000000100000100011100000000000000000000000000000000001100110101010000010101000100100000000000000000010000000000000001100100000000010101010101111011000000000000000000000000000001000") port map( O =>C_28_S_1_L_6_out, I0 =>  inp_feat(82), I1 =>  inp_feat(420), I2 =>  inp_feat(182), I3 =>  inp_feat(451), I4 =>  inp_feat(308), I5 =>  inp_feat(80), I6 =>  inp_feat(339), I7 =>  inp_feat(221)); 
C_28_S_1_L_7_inst : LUT8 generic map(INIT => "0110101010001000000010000000100000000000000000000000000000000000110010100010100000000000000000000000100010000000100110100000100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_1_L_7_out, I0 =>  inp_feat(413), I1 =>  inp_feat(82), I2 =>  inp_feat(144), I3 =>  inp_feat(362), I4 =>  inp_feat(353), I5 =>  inp_feat(148), I6 =>  inp_feat(95), I7 =>  inp_feat(328)); 
C_28_S_2_L_0_inst : LUT8 generic map(INIT => "0011011000001010000000000000010000000000000011000000000000000100110101010000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000010000100000001000000000000000000000000000000000000000000000000") port map( O =>C_28_S_2_L_0_out, I0 =>  inp_feat(81), I1 =>  inp_feat(71), I2 =>  inp_feat(41), I3 =>  inp_feat(247), I4 =>  inp_feat(6), I5 =>  inp_feat(428), I6 =>  inp_feat(238), I7 =>  inp_feat(413)); 
C_28_S_2_L_1_inst : LUT8 generic map(INIT => "0111000001110010000100000100000001010000100000000000000000000000001000100011000000000010000000000010000000000000000000100000000000000000000000001000000000000000010000000000000000100000000000000000000000000000001000000000000000100000000000000000000000000000") port map( O =>C_28_S_2_L_1_out, I0 =>  inp_feat(223), I1 =>  inp_feat(394), I2 =>  inp_feat(331), I3 =>  inp_feat(478), I4 =>  inp_feat(351), I5 =>  inp_feat(303), I6 =>  inp_feat(162), I7 =>  inp_feat(413)); 
C_28_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000100010000000000001011011000010101010100000000000000000000000000010000000100000000000101000001110000000001000000010010001000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_2_L_2_out, I0 =>  inp_feat(158), I1 =>  inp_feat(336), I2 =>  inp_feat(176), I3 =>  inp_feat(164), I4 =>  inp_feat(464), I5 =>  inp_feat(368), I6 =>  inp_feat(30), I7 =>  inp_feat(211)); 
C_28_S_2_L_3_inst : LUT8 generic map(INIT => "0100110001001100010010001100110100000100000001000000000000000001010000000000000000000000000000000000000000000000000000000000000011001100100011000000000000000100110011000000110001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_2_L_3_out, I0 =>  inp_feat(201), I1 =>  inp_feat(98), I2 =>  inp_feat(17), I3 =>  inp_feat(455), I4 =>  inp_feat(478), I5 =>  inp_feat(259), I6 =>  inp_feat(80), I7 =>  inp_feat(339)); 
C_28_S_2_L_4_inst : LUT8 generic map(INIT => "1110000001101100110010101001101010000000010000000001000000000000100010000000101001000000000010010000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000100000000000000000000000") port map( O =>C_28_S_2_L_4_out, I0 =>  inp_feat(382), I1 =>  inp_feat(316), I2 =>  inp_feat(120), I3 =>  inp_feat(30), I4 =>  inp_feat(420), I5 =>  inp_feat(413), I6 =>  inp_feat(95), I7 =>  inp_feat(148)); 
C_28_S_2_L_5_inst : LUT8 generic map(INIT => "0000100000000100010101001000011010001000000000001000100000100000001011000000100001001100100101101000100000000000100010000000000000000000000000000000000000001000100000000000000010001000000000000100000000000100000011000000110010000000000000001000100000000000") port map( O =>C_28_S_2_L_5_out, I0 =>  inp_feat(362), I1 =>  inp_feat(82), I2 =>  inp_feat(52), I3 =>  inp_feat(109), I4 =>  inp_feat(41), I5 =>  inp_feat(18), I6 =>  inp_feat(500), I7 =>  inp_feat(275)); 
C_28_S_2_L_6_inst : LUT8 generic map(INIT => "1010000011100010000000001011000110000000101100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_2_L_6_out, I0 =>  inp_feat(382), I1 =>  inp_feat(420), I2 =>  inp_feat(161), I3 =>  inp_feat(29), I4 =>  inp_feat(500), I5 =>  inp_feat(256), I6 =>  inp_feat(438), I7 =>  inp_feat(282)); 
C_28_S_2_L_7_inst : LUT8 generic map(INIT => "0100011100000010000011100000000000000000000001000000000000011110000010110000010100001101000101110000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000001100001100000001011001010000110100000000000001000000000000000000") port map( O =>C_28_S_2_L_7_out, I0 =>  inp_feat(373), I1 =>  inp_feat(120), I2 =>  inp_feat(221), I3 =>  inp_feat(62), I4 =>  inp_feat(500), I5 =>  inp_feat(148), I6 =>  inp_feat(259), I7 =>  inp_feat(362)); 
C_28_S_3_L_0_inst : LUT8 generic map(INIT => "0100000011000000000000000100010000000000100000000000000010000000000000001000000000000000000000000000000000000000100010001000100011010000100000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_3_L_0_out, I0 =>  inp_feat(37), I1 =>  inp_feat(447), I2 =>  inp_feat(295), I3 =>  inp_feat(31), I4 =>  inp_feat(472), I5 =>  inp_feat(375), I6 =>  inp_feat(304), I7 =>  inp_feat(130)); 
C_28_S_3_L_1_inst : LUT8 generic map(INIT => "1101000111110000100000000000000000010001101000100000000010000000000000000000100000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_3_L_1_out, I0 =>  inp_feat(274), I1 =>  inp_feat(256), I2 =>  inp_feat(328), I3 =>  inp_feat(145), I4 =>  inp_feat(83), I5 =>  inp_feat(480), I6 =>  inp_feat(413), I7 =>  inp_feat(405)); 
C_28_S_3_L_2_inst : LUT8 generic map(INIT => "1111001110100000101000100000000011111011010100110010000000000000010001000100000000000000000000001011001000000011100100000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000001000000100110000") port map( O =>C_28_S_3_L_2_out, I0 =>  inp_feat(336), I1 =>  inp_feat(53), I2 =>  inp_feat(382), I3 =>  inp_feat(82), I4 =>  inp_feat(316), I5 =>  inp_feat(373), I6 =>  inp_feat(141), I7 =>  inp_feat(290)); 
C_28_S_3_L_3_inst : LUT8 generic map(INIT => "0101100000001000110000011000000000000000001000000000000000000000000010101000100011001100101010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_3_L_3_out, I0 =>  inp_feat(177), I1 =>  inp_feat(98), I2 =>  inp_feat(256), I3 =>  inp_feat(262), I4 =>  inp_feat(302), I5 =>  inp_feat(57), I6 =>  inp_feat(244), I7 =>  inp_feat(168)); 
C_28_S_3_L_4_inst : LUT8 generic map(INIT => "0000001000101000001000000000000001010000010100000000000010000000000000001100000000000000000000000000000000000000000000000000000011111000100000000010000000000000000100000101000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_28_S_3_L_4_out, I0 =>  inp_feat(227), I1 =>  inp_feat(265), I2 =>  inp_feat(87), I3 =>  inp_feat(53), I4 =>  inp_feat(313), I5 =>  inp_feat(478), I6 =>  inp_feat(304), I7 =>  inp_feat(460)); 
C_28_S_3_L_5_inst : LUT8 generic map(INIT => "1111001011100011100000000000000000011101001001000000000000000000001000111100001100100001000000000010001010100011000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_3_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(308), I2 =>  inp_feat(239), I3 =>  inp_feat(339), I4 =>  inp_feat(353), I5 =>  inp_feat(420), I6 =>  inp_feat(362), I7 =>  inp_feat(477)); 
C_28_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000100100000000000100010000000000000000000000000000000110000000000000010100000000000000000000000000000000000000000000011001100000000001100101000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_28_S_3_L_6_out, I0 =>  inp_feat(380), I1 =>  inp_feat(98), I2 =>  inp_feat(4), I3 =>  inp_feat(497), I4 =>  inp_feat(86), I5 =>  inp_feat(424), I6 =>  inp_feat(97), I7 =>  inp_feat(75)); 
C_28_S_3_L_7_inst : LUT8 generic map(INIT => "1010101000000000000000001000000000000000000000000000000000000000001100100110101000000000000000000000001100000010000000000000000010011001000000001000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000") port map( O =>C_28_S_3_L_7_out, I0 =>  inp_feat(380), I1 =>  inp_feat(41), I2 =>  inp_feat(256), I3 =>  inp_feat(198), I4 =>  inp_feat(127), I5 =>  inp_feat(372), I6 =>  inp_feat(10), I7 =>  inp_feat(342)); 
C_28_S_4_L_0_inst : LUT8 generic map(INIT => "1110011100001011000000000100011100000000000000000000100000000010000000000000000100000000000000000000000001000000000000000000010000001111110011110000000000001101000000000000000000000010000001100000010100000100000000000000000000001111000001000000110000000000") port map( O =>C_28_S_4_L_0_out, I0 =>  inp_feat(52), I1 =>  inp_feat(327), I2 =>  inp_feat(178), I3 =>  inp_feat(20), I4 =>  inp_feat(351), I5 =>  inp_feat(354), I6 =>  inp_feat(295), I7 =>  inp_feat(259)); 
C_28_S_4_L_1_inst : LUT8 generic map(INIT => "0110101000000001011010100000000000000010000000000010101000000000000000000000000000000000000000001000000010000000101010000010000000000000000000001111000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_4_L_1_out, I0 =>  inp_feat(285), I1 =>  inp_feat(145), I2 =>  inp_feat(238), I3 =>  inp_feat(290), I4 =>  inp_feat(41), I5 =>  inp_feat(468), I6 =>  inp_feat(251), I7 =>  inp_feat(247)); 
C_28_S_4_L_2_inst : LUT8 generic map(INIT => "0000101000000000100111000000000010111000110000001011101000001000110010000000000001011110000010010000100010001000100010100000110100000000000000000000000000000000000100000000000000000000000000000000000000000000000010100000100000000000100000000100001010001000") port map( O =>C_28_S_4_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(420), I2 =>  inp_feat(299), I3 =>  inp_feat(351), I4 =>  inp_feat(259), I5 =>  inp_feat(20), I6 =>  inp_feat(119), I7 =>  inp_feat(182)); 
C_28_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000001010010010001000110001011000000011000000110011001100010010000000101000000000000010000001000000001000000000000000110000000000000000000000000000000000011010100000101000001100000010000010101000101000000010000000001000001000000000000000000000000000") port map( O =>C_28_S_4_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(239), I2 =>  inp_feat(211), I3 =>  inp_feat(97), I4 =>  inp_feat(34), I5 =>  inp_feat(178), I6 =>  inp_feat(227), I7 =>  inp_feat(256)); 
C_28_S_4_L_4_inst : LUT8 generic map(INIT => "1000000100101001010000000000000000010001001100010000000000000000111111110001001000000000000000000000000000010000000000000000000001000000000100000000000000000010000000000000000000000000000000000000000000000010001010100000000000000000000000000000000000000000") port map( O =>C_28_S_4_L_4_out, I0 =>  inp_feat(244), I1 =>  inp_feat(52), I2 =>  inp_feat(20), I3 =>  inp_feat(301), I4 =>  inp_feat(304), I5 =>  inp_feat(445), I6 =>  inp_feat(172), I7 =>  inp_feat(380)); 
C_28_S_4_L_5_inst : LUT8 generic map(INIT => "0000100000001110000100000000000011001100000000100000000000000000000000000000000000000000000000000000000000010100000000000000000001011100000000000011000000000000110011000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000") port map( O =>C_28_S_4_L_5_out, I0 =>  inp_feat(308), I1 =>  inp_feat(407), I2 =>  inp_feat(256), I3 =>  inp_feat(105), I4 =>  inp_feat(251), I5 =>  inp_feat(300), I6 =>  inp_feat(80), I7 =>  inp_feat(339)); 
C_28_S_4_L_6_inst : LUT8 generic map(INIT => "1111000000110010001100001011000010110000000010001111000000101000000000000000000000000000000000000000000000101000000000100000001000000010100000000000001001100000000010000000000000100000001010000000000000000000000010000000000000000010000000000000101000001000") port map( O =>C_28_S_4_L_6_out, I0 =>  inp_feat(93), I1 =>  inp_feat(299), I2 =>  inp_feat(354), I3 =>  inp_feat(120), I4 =>  inp_feat(201), I5 =>  inp_feat(19), I6 =>  inp_feat(182), I7 =>  inp_feat(164)); 
C_28_S_4_L_7_inst : LUT8 generic map(INIT => "0000010011000000010000000100000010000000100010000001010000001000000000000000000000000000000000000000001000000000000000000000001001000000110000001000101011000000000000001100000011000101110000000000000000000000000000000000000000000000000000000000100000000000") port map( O =>C_28_S_4_L_7_out, I0 =>  inp_feat(20), I1 =>  inp_feat(295), I2 =>  inp_feat(286), I3 =>  inp_feat(93), I4 =>  inp_feat(177), I5 =>  inp_feat(238), I6 =>  inp_feat(80), I7 =>  inp_feat(339)); 
C_29_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000000010000100000000101100000010000000100000000000000010000000100000100000000000000000000000000000000000110000000000001011000000000000101101000001000000000000000000100000000000000010100000000000001010000000000000") port map( O =>C_29_S_0_L_0_out, I0 =>  inp_feat(362), I1 =>  inp_feat(130), I2 =>  inp_feat(371), I3 =>  inp_feat(161), I4 =>  inp_feat(20), I5 =>  inp_feat(221), I6 =>  inp_feat(211), I7 =>  inp_feat(299)); 
C_29_S_0_L_1_inst : LUT8 generic map(INIT => "1000000000000000000000000000000000000000000000000000000000000000100010001000000000101010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_0_L_1_out, I0 =>  inp_feat(126), I1 =>  inp_feat(504), I2 =>  inp_feat(412), I3 =>  inp_feat(506), I4 =>  inp_feat(82), I5 =>  inp_feat(424), I6 =>  inp_feat(223), I7 =>  inp_feat(83)); 
C_29_S_0_L_2_inst : LUT8 generic map(INIT => "0111010100000000010100000000000010100010000000000000000000000000000000000000000000000000000000000000100000000010000000000000000011110000000000000000000000000000111100000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000") port map( O =>C_29_S_0_L_2_out, I0 =>  inp_feat(144), I1 =>  inp_feat(201), I2 =>  inp_feat(336), I3 =>  inp_feat(98), I4 =>  inp_feat(30), I5 =>  inp_feat(121), I6 =>  inp_feat(13), I7 =>  inp_feat(223)); 
C_29_S_0_L_3_inst : LUT8 generic map(INIT => "0000101000000000000010000000100011001100000011000000110000001100000000000000000000000000000010000000000000000000000010000000100010001000100000001000100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_0_L_3_out, I0 =>  inp_feat(161), I1 =>  inp_feat(290), I2 =>  inp_feat(221), I3 =>  inp_feat(331), I4 =>  inp_feat(339), I5 =>  inp_feat(41), I6 =>  inp_feat(354), I7 =>  inp_feat(25)); 
C_29_S_0_L_4_inst : LUT8 generic map(INIT => "0000000100000010000100000001000011110001100000000000000000000000000000000000000000000000000000000000000000000000010000000000000011010000011111100000000000000000101100001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_0_L_4_out, I0 =>  inp_feat(387), I1 =>  inp_feat(29), I2 =>  inp_feat(40), I3 =>  inp_feat(97), I4 =>  inp_feat(408), I5 =>  inp_feat(300), I6 =>  inp_feat(477), I7 =>  inp_feat(17)); 
C_29_S_0_L_5_inst : LUT8 generic map(INIT => "1100100010000000100000001000101000000000000000001000000010001000000000000000000000000000000010000000000000000000000000000000100000000000000000001000000000000000000000000000000010110000100010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_0_L_5_out, I0 =>  inp_feat(98), I1 =>  inp_feat(336), I2 =>  inp_feat(58), I3 =>  inp_feat(308), I4 =>  inp_feat(29), I5 =>  inp_feat(186), I6 =>  inp_feat(304), I7 =>  inp_feat(161)); 
C_29_S_0_L_6_inst : LUT8 generic map(INIT => "0000000010000000110100000000010000000000000000000000000100000100000000000000000001000000000000000000000000000000000000000000000011000000110001000000000000001100001000001000110011000000000000001000000001000000000001000000000000000000000000000000000000000100") port map( O =>C_29_S_0_L_6_out, I0 =>  inp_feat(52), I1 =>  inp_feat(183), I2 =>  inp_feat(362), I3 =>  inp_feat(144), I4 =>  inp_feat(220), I5 =>  inp_feat(354), I6 =>  inp_feat(316), I7 =>  inp_feat(299)); 
C_29_S_0_L_7_inst : LUT8 generic map(INIT => "0101001000010010000010100010001000100010001000000000000000000010001010100110001000100010111000100000100000000000000000000111001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_0_L_7_out, I0 =>  inp_feat(158), I1 =>  inp_feat(221), I2 =>  inp_feat(17), I3 =>  inp_feat(340), I4 =>  inp_feat(399), I5 =>  inp_feat(273), I6 =>  inp_feat(509), I7 =>  inp_feat(64)); 
C_29_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000000010000100000000101100000010000000100000000000000010000000100000100000000000000000000000000000000000110000000000001011000000000000101101000001000000000000000000100000000000000010100000000000001010000000000000") port map( O =>C_29_S_1_L_0_out, I0 =>  inp_feat(362), I1 =>  inp_feat(130), I2 =>  inp_feat(371), I3 =>  inp_feat(161), I4 =>  inp_feat(20), I5 =>  inp_feat(221), I6 =>  inp_feat(211), I7 =>  inp_feat(299)); 
C_29_S_1_L_1_inst : LUT8 generic map(INIT => "1111110100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_1_L_1_out, I0 =>  inp_feat(37), I1 =>  inp_feat(94), I2 =>  inp_feat(407), I3 =>  inp_feat(355), I4 =>  inp_feat(69), I5 =>  inp_feat(370), I6 =>  inp_feat(353), I7 =>  inp_feat(506)); 
C_29_S_1_L_2_inst : LUT8 generic map(INIT => "1101000000100000111110001000100000000000000000000100000000001000000100000000000010000000000000100000000000000000000000000000000000100000000000000010000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000") port map( O =>C_29_S_1_L_2_out, I0 =>  inp_feat(464), I1 =>  inp_feat(339), I2 =>  inp_feat(158), I3 =>  inp_feat(336), I4 =>  inp_feat(201), I5 =>  inp_feat(98), I6 =>  inp_feat(354), I7 =>  inp_feat(30)); 
C_29_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000001000000000000000101000000000000000000000000000000000000000000000101000001000000000000000000010101000100000001000100010000000100010000000000010001000100000000000000000000000100000000000000000000000000000001000000000000000") port map( O =>C_29_S_1_L_3_out, I0 =>  inp_feat(331), I1 =>  inp_feat(4), I2 =>  inp_feat(229), I3 =>  inp_feat(445), I4 =>  inp_feat(117), I5 =>  inp_feat(256), I6 =>  inp_feat(378), I7 =>  inp_feat(223)); 
C_29_S_1_L_4_inst : LUT8 generic map(INIT => "0000001100001101001000000000000000000000000001001000100000000010010010000000001010001010100010100000000000001000001010100000101000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_1_L_4_out, I0 =>  inp_feat(86), I1 =>  inp_feat(430), I2 =>  inp_feat(29), I3 =>  inp_feat(346), I4 =>  inp_feat(178), I5 =>  inp_feat(308), I6 =>  inp_feat(464), I7 =>  inp_feat(492)); 
C_29_S_1_L_5_inst : LUT8 generic map(INIT => "1010000000000000001000000000000010100010000000000000000000000000000000000000101000000000000000000000000000000000000000000000000011000000000000001010000000000000101000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_1_L_5_out, I0 =>  inp_feat(217), I1 =>  inp_feat(52), I2 =>  inp_feat(162), I3 =>  inp_feat(390), I4 =>  inp_feat(493), I5 =>  inp_feat(244), I6 =>  inp_feat(304), I7 =>  inp_feat(265)); 
C_29_S_1_L_6_inst : LUT8 generic map(INIT => "1100010000000000010011000000010000000000000000000000010000000000100000010000000011001101000000000000000000000000000000001000000001001000000000001101110000010000000000000000000011000000000000000000100000000000110011000000000000000000000000000000000000000000") port map( O =>C_29_S_1_L_6_out, I0 =>  inp_feat(41), I1 =>  inp_feat(468), I2 =>  inp_feat(399), I3 =>  inp_feat(344), I4 =>  inp_feat(302), I5 =>  inp_feat(322), I6 =>  inp_feat(244), I7 =>  inp_feat(144)); 
C_29_S_1_L_7_inst : LUT8 generic map(INIT => "0100010001001000000100010000000001000000110000000100001011000100000000000000000000000001000000000000000000000000000000000000000001000100110011000101000111001100010000111100110000000111110011000000000000000000000001000000000000000000000000000000000100000000") port map( O =>C_29_S_1_L_7_out, I0 =>  inp_feat(144), I1 =>  inp_feat(331), I2 =>  inp_feat(238), I3 =>  inp_feat(93), I4 =>  inp_feat(241), I5 =>  inp_feat(222), I6 =>  inp_feat(161), I7 =>  inp_feat(339)); 
C_29_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000000010000100000000101100000010000000100000000000000010000000100000100000000000000000000000000000000000110000000000001011000000000000101101000001000000000000000000100000000000000010100000000000001010000000000000") port map( O =>C_29_S_2_L_0_out, I0 =>  inp_feat(362), I1 =>  inp_feat(130), I2 =>  inp_feat(371), I3 =>  inp_feat(161), I4 =>  inp_feat(20), I5 =>  inp_feat(221), I6 =>  inp_feat(211), I7 =>  inp_feat(299)); 
C_29_S_2_L_1_inst : LUT8 generic map(INIT => "1011001011000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_2_L_1_out, I0 =>  inp_feat(189), I1 =>  inp_feat(108), I2 =>  inp_feat(55), I3 =>  inp_feat(199), I4 =>  inp_feat(355), I5 =>  inp_feat(370), I6 =>  inp_feat(353), I7 =>  inp_feat(506)); 
C_29_S_2_L_2_inst : LUT8 generic map(INIT => "1111000000100001101000000000000001110000011111111010000011100000000000000000000000000000000000000000000001000010000000000000000000000000000000010000000010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_2_L_2_out, I0 =>  inp_feat(484), I1 =>  inp_feat(37), I2 =>  inp_feat(158), I3 =>  inp_feat(201), I4 =>  inp_feat(144), I5 =>  inp_feat(509), I6 =>  inp_feat(98), I7 =>  inp_feat(38)); 
C_29_S_2_L_3_inst : LUT8 generic map(INIT => "0010000000000000000000000010000110000000000000000010000000000000000000000000000000000000000000000000000000000000001101100000000010100000000000000010000010010000101000000000000010100000000000000000000000000000001000000000000000100000000000000000000000000000") port map( O =>C_29_S_2_L_3_out, I0 =>  inp_feat(309), I1 =>  inp_feat(244), I2 =>  inp_feat(98), I3 =>  inp_feat(64), I4 =>  inp_feat(478), I5 =>  inp_feat(256), I6 =>  inp_feat(378), I7 =>  inp_feat(223)); 
C_29_S_2_L_4_inst : LUT8 generic map(INIT => "0100001100000001101010100000000000011001001000010000000000000100000000000000000000000000000000000000000000000000000000000000000011100000000000001010101000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000") port map( O =>C_29_S_2_L_4_out, I0 =>  inp_feat(318), I1 =>  inp_feat(256), I2 =>  inp_feat(244), I3 =>  inp_feat(492), I4 =>  inp_feat(17), I5 =>  inp_feat(7), I6 =>  inp_feat(344), I7 =>  inp_feat(394)); 
C_29_S_2_L_5_inst : LUT8 generic map(INIT => "1100100011000000110001001100010000000000000001010000010001000100000000001100000011000000110000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_2_L_5_out, I0 =>  inp_feat(308), I1 =>  inp_feat(161), I2 =>  inp_feat(331), I3 =>  inp_feat(144), I4 =>  inp_feat(339), I5 =>  inp_feat(30), I6 =>  inp_feat(346), I7 =>  inp_feat(336)); 
C_29_S_2_L_6_inst : LUT8 generic map(INIT => "0101100101010000000000000000110011100100111110000000000010000100000000000000000000000000000000001100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_29_S_2_L_6_out, I0 =>  inp_feat(244), I1 =>  inp_feat(233), I2 =>  inp_feat(445), I3 =>  inp_feat(12), I4 =>  inp_feat(64), I5 =>  inp_feat(223), I6 =>  inp_feat(74), I7 =>  inp_feat(474)); 
C_29_S_2_L_7_inst : LUT8 generic map(INIT => "0000000010000000100001000000000000000000000000000000000000000000100000000100000000000000010000000000000000000000000000000000000010101000111010001000000011000100000000000000001000000010010000000000000010000100000000000100000000000000000000000000000000000000") port map( O =>C_29_S_2_L_7_out, I0 =>  inp_feat(247), I1 =>  inp_feat(472), I2 =>  inp_feat(431), I3 =>  inp_feat(256), I4 =>  inp_feat(265), I5 =>  inp_feat(290), I6 =>  inp_feat(465), I7 =>  inp_feat(75)); 
C_29_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000000010000100000000101100000010000000100000000000000010000000100000100000000000000000000000000000000000110000000000001011000000000000101101000001000000000000000000100000000000000010100000000000001010000000000000") port map( O =>C_29_S_3_L_0_out, I0 =>  inp_feat(362), I1 =>  inp_feat(130), I2 =>  inp_feat(371), I3 =>  inp_feat(161), I4 =>  inp_feat(20), I5 =>  inp_feat(221), I6 =>  inp_feat(211), I7 =>  inp_feat(299)); 
C_29_S_3_L_1_inst : LUT8 generic map(INIT => "1011001011000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_3_L_1_out, I0 =>  inp_feat(189), I1 =>  inp_feat(108), I2 =>  inp_feat(55), I3 =>  inp_feat(199), I4 =>  inp_feat(370), I5 =>  inp_feat(355), I6 =>  inp_feat(353), I7 =>  inp_feat(506)); 
C_29_S_3_L_2_inst : LUT8 generic map(INIT => "1111000000100001101000000000000001110000011111111010000011100000000000000000000000000000000000000000000001000010000000000000000000000000000000010000000010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_3_L_2_out, I0 =>  inp_feat(484), I1 =>  inp_feat(37), I2 =>  inp_feat(158), I3 =>  inp_feat(201), I4 =>  inp_feat(144), I5 =>  inp_feat(509), I6 =>  inp_feat(98), I7 =>  inp_feat(38)); 
C_29_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000011000000010010000000000000000000001000000000000000000000000000000001000000000000000000000000001100100001000011010100000011000000010000001001110011000000000000000100100000000000000000000000000010000000000000001000000000000000000000000000") port map( O =>C_29_S_3_L_3_out, I0 =>  inp_feat(97), I1 =>  inp_feat(435), I2 =>  inp_feat(134), I3 =>  inp_feat(445), I4 =>  inp_feat(478), I5 =>  inp_feat(256), I6 =>  inp_feat(378), I7 =>  inp_feat(223)); 
C_29_S_3_L_4_inst : LUT8 generic map(INIT => "0000000011100000110010000110000000000000000000000000000000000000010000001100000011000000111000000000000000000000000000000000000000000000100000000000000001000000010000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000") port map( O =>C_29_S_3_L_4_out, I0 =>  inp_feat(94), I1 =>  inp_feat(324), I2 =>  inp_feat(304), I3 =>  inp_feat(223), I4 =>  inp_feat(373), I5 =>  inp_feat(336), I6 =>  inp_feat(300), I7 =>  inp_feat(478)); 
C_29_S_3_L_5_inst : LUT8 generic map(INIT => "0101110000010001000001110001011000000000000000000000000000000000110010010000010000000000000000000000000000000000000000000000000011110000111101110000000000000100001000000000000000000000000000001111100011111111000000000000000000000000000000000000000000000000") port map( O =>C_29_S_3_L_5_out, I0 =>  inp_feat(144), I1 =>  inp_feat(367), I2 =>  inp_feat(238), I3 =>  inp_feat(339), I4 =>  inp_feat(30), I5 =>  inp_feat(307), I6 =>  inp_feat(300), I7 =>  inp_feat(464)); 
C_29_S_3_L_6_inst : LUT8 generic map(INIT => "0010000000100000101000101010000000100000001010000010100000100000000000000000000000000000000000000000000001000000000000000000000010100000101110001010000000110000001000001011000000000000101000110000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_29_S_3_L_6_out, I0 =>  inp_feat(336), I1 =>  inp_feat(130), I2 =>  inp_feat(199), I3 =>  inp_feat(340), I4 =>  inp_feat(505), I5 =>  inp_feat(430), I6 =>  inp_feat(322), I7 =>  inp_feat(244)); 
C_29_S_3_L_7_inst : LUT8 generic map(INIT => "0010010010110010101000000000000000000000000000000000000000000000101110000000000011110000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_29_S_3_L_7_out, I0 =>  inp_feat(316), I1 =>  inp_feat(339), I2 =>  inp_feat(183), I3 =>  inp_feat(331), I4 =>  inp_feat(97), I5 =>  inp_feat(403), I6 =>  inp_feat(15), I7 =>  inp_feat(344)); 
C_29_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000000010000100000000101100000010000000100000000000000010000000100000100000000000000000000000000000000000110000000000001011000000000000101101000001000000000000000000100000000000000010100000000000001010000000000000") port map( O =>C_29_S_4_L_0_out, I0 =>  inp_feat(362), I1 =>  inp_feat(130), I2 =>  inp_feat(371), I3 =>  inp_feat(161), I4 =>  inp_feat(20), I5 =>  inp_feat(221), I6 =>  inp_feat(211), I7 =>  inp_feat(299)); 
C_29_S_4_L_1_inst : LUT8 generic map(INIT => "1110101011100000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000010000000100000000000000000000000000000000000000000") port map( O =>C_29_S_4_L_1_out, I0 =>  inp_feat(331), I1 =>  inp_feat(130), I2 =>  inp_feat(324), I3 =>  inp_feat(380), I4 =>  inp_feat(370), I5 =>  inp_feat(353), I6 =>  inp_feat(355), I7 =>  inp_feat(506)); 
C_29_S_4_L_2_inst : LUT8 generic map(INIT => "1110111000101110000000000100100011101010000010000000100000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_4_L_2_out, I0 =>  inp_feat(328), I1 =>  inp_feat(144), I2 =>  inp_feat(464), I3 =>  inp_feat(58), I4 =>  inp_feat(431), I5 =>  inp_feat(37), I6 =>  inp_feat(331), I7 =>  inp_feat(385)); 
C_29_S_4_L_3_inst : LUT8 generic map(INIT => "0000111000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101010000000001000000000000000101000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_4_L_3_out, I0 =>  inp_feat(53), I1 =>  inp_feat(308), I2 =>  inp_feat(144), I3 =>  inp_feat(161), I4 =>  inp_feat(328), I5 =>  inp_feat(286), I6 =>  inp_feat(477), I7 =>  inp_feat(464)); 
C_29_S_4_L_4_inst : LUT8 generic map(INIT => "0010000010100000000000000000001100101000001100110000000000000000100000001000000000000000000000000000000000000000000000000000000010100000101000100000000010100010000000000010000000010001000011000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_4_L_4_out, I0 =>  inp_feat(7), I1 =>  inp_feat(157), I2 =>  inp_feat(239), I3 =>  inp_feat(244), I4 =>  inp_feat(247), I5 =>  inp_feat(372), I6 =>  inp_feat(263), I7 =>  inp_feat(256)); 
C_29_S_4_L_5_inst : LUT8 generic map(INIT => "0100110111000000000000000000000011001010000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_29_S_4_L_5_out, I0 =>  inp_feat(144), I1 =>  inp_feat(82), I2 =>  inp_feat(31), I3 =>  inp_feat(304), I4 =>  inp_feat(247), I5 =>  inp_feat(18), I6 =>  inp_feat(306), I7 =>  inp_feat(478)); 
C_29_S_4_L_6_inst : LUT8 generic map(INIT => "1010010000001000100010000000000010001100000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000010000000000000000000000000000000000000000001000100000000000000000000000000") port map( O =>C_29_S_4_L_6_out, I0 =>  inp_feat(45), I1 =>  inp_feat(36), I2 =>  inp_feat(256), I3 =>  inp_feat(231), I4 =>  inp_feat(346), I5 =>  inp_feat(37), I6 =>  inp_feat(295), I7 =>  inp_feat(224)); 
C_29_S_4_L_7_inst : LUT8 generic map(INIT => "0111000010000000111100000000000001110000000000000111001100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010100000000000000000000000000000") port map( O =>C_29_S_4_L_7_out, I0 =>  inp_feat(157), I1 =>  inp_feat(256), I2 =>  inp_feat(98), I3 =>  inp_feat(283), I4 =>  inp_feat(346), I5 =>  inp_feat(37), I6 =>  inp_feat(80), I7 =>  inp_feat(290)); 
C_30_S_0_L_0_inst : LUT8 generic map(INIT => "0101000000000000000000000000000011000000110000001101000000000100000000000000000000000000000000001000001000000000100000000000000010000000000000001010000000000000110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_0_L_0_out, I0 =>  inp_feat(388), I1 =>  inp_feat(183), I2 =>  inp_feat(258), I3 =>  inp_feat(435), I4 =>  inp_feat(331), I5 =>  inp_feat(464), I6 =>  inp_feat(474), I7 =>  inp_feat(299)); 
C_30_S_0_L_1_inst : LUT8 generic map(INIT => "0000010000001000000000000000110111001100000011000100000000000000000000000000000000000001000001110000000000000000000000000000000010100000100010001110000010001000110011001100100011000000110000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_0_L_1_out, I0 =>  inp_feat(93), I1 =>  inp_feat(331), I2 =>  inp_feat(452), I3 =>  inp_feat(77), I4 =>  inp_feat(95), I5 =>  inp_feat(223), I6 =>  inp_feat(421), I7 =>  inp_feat(29)); 
C_30_S_0_L_2_inst : LUT8 generic map(INIT => "1010000010000000000000000000000010000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010101000100000100000000000000000111100001010000001000100001000000000000000000000000000000000000010100000111000000100000010000000") port map( O =>C_30_S_0_L_2_out, I0 =>  inp_feat(306), I1 =>  inp_feat(493), I2 =>  inp_feat(472), I3 =>  inp_feat(40), I4 =>  inp_feat(57), I5 =>  inp_feat(195), I6 =>  inp_feat(100), I7 =>  inp_feat(41)); 
C_30_S_0_L_3_inst : LUT8 generic map(INIT => "0010111101100010000000100000000000001111000001000010001000000010110011100000101000000000000000000000001000000100000000000000000011111111000000000000000000000000011001100010000000100010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_0_L_3_out, I0 =>  inp_feat(20), I1 =>  inp_feat(201), I2 =>  inp_feat(373), I3 =>  inp_feat(413), I4 =>  inp_feat(148), I5 =>  inp_feat(182), I6 =>  inp_feat(247), I7 =>  inp_feat(144)); 
C_30_S_0_L_4_inst : LUT8 generic map(INIT => "1010110001101100000010000000100011110001101010100000000000000000101000000000000000000000000000001011000000000000000010000000000000000100000000000000100000000000101010000000001000000000000000000000000000000000100001000000000000000000000000000000000000000000") port map( O =>C_30_S_0_L_4_out, I0 =>  inp_feat(183), I1 =>  inp_feat(222), I2 =>  inp_feat(31), I3 =>  inp_feat(351), I4 =>  inp_feat(167), I5 =>  inp_feat(509), I6 =>  inp_feat(7), I7 =>  inp_feat(413)); 
C_30_S_0_L_5_inst : LUT8 generic map(INIT => "1110100000000101000000000000000010110000010100010010000000000000110011000000000000000000000000001000101000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_0_L_5_out, I0 =>  inp_feat(41), I1 =>  inp_feat(478), I2 =>  inp_feat(476), I3 =>  inp_feat(492), I4 =>  inp_feat(490), I5 =>  inp_feat(61), I6 =>  inp_feat(18), I7 =>  inp_feat(405)); 
C_30_S_0_L_6_inst : LUT8 generic map(INIT => "0010001000101010001000101010000000000000000000000000000000000000100010001010100011000000101000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001010100000000000000000000000000000000000") port map( O =>C_30_S_0_L_6_out, I0 =>  inp_feat(504), I1 =>  inp_feat(300), I2 =>  inp_feat(102), I3 =>  inp_feat(312), I4 =>  inp_feat(256), I5 =>  inp_feat(140), I6 =>  inp_feat(448), I7 =>  inp_feat(143)); 
C_30_S_0_L_7_inst : LUT8 generic map(INIT => "1000000010001010100010000001000100000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000010111010110000101100110011111000000010000000000001000100000000000101100010000000000000001110100000000000000000000000000000000000") port map( O =>C_30_S_0_L_7_out, I0 =>  inp_feat(82), I1 =>  inp_feat(290), I2 =>  inp_feat(420), I3 =>  inp_feat(158), I4 =>  inp_feat(221), I5 =>  inp_feat(247), I6 =>  inp_feat(353), I7 =>  inp_feat(178)); 
C_30_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000100000001001000000000000000000000000000101000100010000101000000000000010100000000000000000000000000000000000000000000010110000001100001010001000010000000000000000000000000000000000000010000000000000101000000000000000000000000000000000000000000000") port map( O =>C_30_S_1_L_0_out, I0 =>  inp_feat(492), I1 =>  inp_feat(291), I2 =>  inp_feat(57), I3 =>  inp_feat(36), I4 =>  inp_feat(29), I5 =>  inp_feat(100), I6 =>  inp_feat(34), I7 =>  inp_feat(75)); 
C_30_S_1_L_1_inst : LUT8 generic map(INIT => "0001000001000100100000001101010100010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000011010000110100011000000011000001000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_1_L_1_out, I0 =>  inp_feat(509), I1 =>  inp_feat(376), I2 =>  inp_feat(310), I3 =>  inp_feat(29), I4 =>  inp_feat(256), I5 =>  inp_feat(57), I6 =>  inp_feat(438), I7 =>  inp_feat(157)); 
C_30_S_1_L_2_inst : LUT8 generic map(INIT => "1110100000000000100000000010000010000000000000000000100000000000101111110000010010100000100000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000010000000000000000000000001000000000000000000000000") port map( O =>C_30_S_1_L_2_out, I0 =>  inp_feat(6), I1 =>  inp_feat(265), I2 =>  inp_feat(492), I3 =>  inp_feat(57), I4 =>  inp_feat(472), I5 =>  inp_feat(36), I6 =>  inp_feat(29), I7 =>  inp_feat(100)); 
C_30_S_1_L_3_inst : LUT8 generic map(INIT => "1101010101010001000001000000000010000010000100010000000010000000000000000100000000000000000000000000100000000000000000000000000011111010111100000000000010000000101000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_1_L_3_out, I0 =>  inp_feat(509), I1 =>  inp_feat(256), I2 =>  inp_feat(247), I3 =>  inp_feat(457), I4 =>  inp_feat(331), I5 =>  inp_feat(342), I6 =>  inp_feat(490), I7 =>  inp_feat(18)); 
C_30_S_1_L_4_inst : LUT8 generic map(INIT => "1000000010110010110000000000000000000000010000000100000000100000100000001110000100100000000000000001000000100000000000000010000011000000100010010000000000000000000000000010000000000000001000000000000010001000000000000000100011100000111000100000000000100010") port map( O =>C_30_S_1_L_4_out, I0 =>  inp_feat(468), I1 =>  inp_feat(372), I2 =>  inp_feat(98), I3 =>  inp_feat(77), I4 =>  inp_feat(153), I5 =>  inp_feat(38), I6 =>  inp_feat(484), I7 =>  inp_feat(275)); 
C_30_S_1_L_5_inst : LUT8 generic map(INIT => "0011000110010001000100010001100100000000000000000000010000000000001000001001000001000000111000100000000000000000000000000000000000011100110111000101000001010000000000001100000001000000010100000100001000000010000000001100000000000000000000000000000000000000") port map( O =>C_30_S_1_L_5_out, I0 =>  inp_feat(178), I1 =>  inp_feat(303), I2 =>  inp_feat(290), I3 =>  inp_feat(201), I4 =>  inp_feat(373), I5 =>  inp_feat(477), I6 =>  inp_feat(420), I7 =>  inp_feat(458)); 
C_30_S_1_L_6_inst : LUT8 generic map(INIT => "0101000011000000111100000000000000000000000000001101000000000000010100000000000011010000001000100101000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_30_S_1_L_6_out, I0 =>  inp_feat(75), I1 =>  inp_feat(265), I2 =>  inp_feat(79), I3 =>  inp_feat(143), I4 =>  inp_feat(29), I5 =>  inp_feat(124), I6 =>  inp_feat(434), I7 =>  inp_feat(405)); 
C_30_S_1_L_7_inst : LUT8 generic map(INIT => "0100100000000000000000000000000000000001111001000000000000000000001000001101100100000000000000000000001010100000001000000000000010101000000000000000000000000000000000000000000000100000001000001010000000000000100000000000000000000000000000000000000000000000") port map( O =>C_30_S_1_L_7_out, I0 =>  inp_feat(331), I1 =>  inp_feat(373), I2 =>  inp_feat(504), I3 =>  inp_feat(351), I4 =>  inp_feat(96), I5 =>  inp_feat(87), I6 =>  inp_feat(365), I7 =>  inp_feat(433)); 
C_30_S_2_L_0_inst : LUT8 generic map(INIT => "0010111000010010100011000000000000000000000001000000000000000000000000101000001000100101000000000000000000000000000000000000000000000100110011101100100010101011000000000000101000000000100010000000000100010000000000001000100000000000000000000000000000000000") port map( O =>C_30_S_2_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(53), I2 =>  inp_feat(52), I3 =>  inp_feat(449), I4 =>  inp_feat(95), I5 =>  inp_feat(353), I6 =>  inp_feat(413), I7 =>  inp_feat(241)); 
C_30_S_2_L_1_inst : LUT8 generic map(INIT => "1101011001000001000101000001000011100100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000011011101000001011110000000000000000000000000010000000000000000000000000101000101000000000000000000000000000000000000000000000000") port map( O =>C_30_S_2_L_1_out, I0 =>  inp_feat(99), I1 =>  inp_feat(493), I2 =>  inp_feat(411), I3 =>  inp_feat(492), I4 =>  inp_feat(472), I5 =>  inp_feat(36), I6 =>  inp_feat(100), I7 =>  inp_feat(29)); 
C_30_S_2_L_2_inst : LUT8 generic map(INIT => "1001011000000100000010010000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101000000001001100000010000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_2_L_2_out, I0 =>  inp_feat(391), I1 =>  inp_feat(364), I2 =>  inp_feat(228), I3 =>  inp_feat(328), I4 =>  inp_feat(186), I5 =>  inp_feat(112), I6 =>  inp_feat(140), I7 =>  inp_feat(434)); 
C_30_S_2_L_3_inst : LUT8 generic map(INIT => "0010000000000010111000001000000000000000000000000000000010000000110000000000000010000000000000000000000000000000000000000000000010110010001000000111000010110000000000100000000001000000000000001000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_30_S_2_L_3_out, I0 =>  inp_feat(290), I1 =>  inp_feat(51), I2 =>  inp_feat(182), I3 =>  inp_feat(6), I4 =>  inp_feat(434), I5 =>  inp_feat(148), I6 =>  inp_feat(18), I7 =>  inp_feat(166)); 
C_30_S_2_L_4_inst : LUT8 generic map(INIT => "1001010100000101110001010000000100000100000000000000010000000001011111111001101110000000000000000000111100000000000010000000000011000110000000000100010000000000010011000000100010001100000000000100111000000010100010100000101000001110000000000000000000000000") port map( O =>C_30_S_2_L_4_out, I0 =>  inp_feat(228), I1 =>  inp_feat(238), I2 =>  inp_feat(75), I3 =>  inp_feat(416), I4 =>  inp_feat(53), I5 =>  inp_feat(256), I6 =>  inp_feat(277), I7 =>  inp_feat(77)); 
C_30_S_2_L_5_inst : LUT8 generic map(INIT => "0010111000001000100111100100000000000010000000000000000011000000000000100000100000000000000000000000001000000000000000000000000000000000000000000111110001000000000000000100000011100000010000000000000001000000010000001100000000000000000000000000000001000000") port map( O =>C_30_S_2_L_5_out, I0 =>  inp_feat(222), I1 =>  inp_feat(102), I2 =>  inp_feat(223), I3 =>  inp_feat(176), I4 =>  inp_feat(494), I5 =>  inp_feat(413), I6 =>  inp_feat(374), I7 =>  inp_feat(308)); 
C_30_S_2_L_6_inst : LUT8 generic map(INIT => "0000110000100000001000001100000011100100000000001110110000001000010000000000000010000100000000100000000000000000000011000000000011010100110000000000000000000000000000000000000000000000000000000010000000110010000000000000000011000100000000000000000000000100") port map( O =>C_30_S_2_L_6_out, I0 =>  inp_feat(115), I1 =>  inp_feat(218), I2 =>  inp_feat(141), I3 =>  inp_feat(413), I4 =>  inp_feat(95), I5 =>  inp_feat(144), I6 =>  inp_feat(480), I7 =>  inp_feat(74)); 
C_30_S_2_L_7_inst : LUT8 generic map(INIT => "1001000001000000000000100000000010000000110000000000000000000000000000101011100000000000000100001101111111010000110000001100011011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000") port map( O =>C_30_S_2_L_7_out, I0 =>  inp_feat(238), I1 =>  inp_feat(477), I2 =>  inp_feat(331), I3 =>  inp_feat(18), I4 =>  inp_feat(98), I5 =>  inp_feat(77), I6 =>  inp_feat(105), I7 =>  inp_feat(184)); 
C_30_S_3_L_0_inst : LUT8 generic map(INIT => "0000000010000000011000000000000000100000000000001110000000000000000000001000000010011000110000000010101000000000111111010000101100000000000000001000000000000000000000000000000000000000000000001000100000000000100000000000000010100000000000001010000000000000") port map( O =>C_30_S_3_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(73), I2 =>  inp_feat(60), I3 =>  inp_feat(506), I4 =>  inp_feat(29), I5 =>  inp_feat(256), I6 =>  inp_feat(434), I7 =>  inp_feat(124)); 
C_30_S_3_L_1_inst : LUT8 generic map(INIT => "0010000000000010000000000000000000101000000000000000000000000000001010000000000010000000000000001010101100000000000000000000000010101000100000100000000000000000101010000000000000000000000000001010000010001010000000001000101010100000000000000000000000000000") port map( O =>C_30_S_3_L_1_out, I0 =>  inp_feat(57), I1 =>  inp_feat(37), I2 =>  inp_feat(53), I3 =>  inp_feat(501), I4 =>  inp_feat(237), I5 =>  inp_feat(256), I6 =>  inp_feat(77), I7 =>  inp_feat(277)); 
C_30_S_3_L_2_inst : LUT8 generic map(INIT => "0000100000000001000000100000001000000000000000000000000000000000101010100000100000111000001000001000010000000000100010000000000010001010000000000000001000000000000000000000000000000000000000000100100010001010000000101010101011001101000010001000110000101010") port map( O =>C_30_S_3_L_2_out, I0 =>  inp_feat(477), I1 =>  inp_feat(316), I2 =>  inp_feat(52), I3 =>  inp_feat(331), I4 =>  inp_feat(420), I5 =>  inp_feat(182), I6 =>  inp_feat(71), I7 =>  inp_feat(210)); 
C_30_S_3_L_3_inst : LUT8 generic map(INIT => "0010110010101000111000110110110011110010001000011110000111101010000000001000000011000000000000000100000001000000000000000100000000010000000000000000000010000000000000000000000000000000000000001101000010000000100000000000000000000000000000000000000000000000") port map( O =>C_30_S_3_L_3_out, I0 =>  inp_feat(53), I1 =>  inp_feat(18), I2 =>  inp_feat(427), I3 =>  inp_feat(120), I4 =>  inp_feat(238), I5 =>  inp_feat(259), I6 =>  inp_feat(74), I7 =>  inp_feat(131)); 
C_30_S_3_L_4_inst : LUT8 generic map(INIT => "1000000000000010100000000000000010000000010000001000000000000000100000011010000010000000000000001000100011100000000001001100000000000000000000000000000000000000000000000000000000000000000000000000000001000011010000000110100000000000110000000000000000000000") port map( O =>C_30_S_3_L_4_out, I0 =>  inp_feat(6), I1 =>  inp_feat(306), I2 =>  inp_feat(57), I3 =>  inp_feat(174), I4 =>  inp_feat(40), I5 =>  inp_feat(493), I6 =>  inp_feat(29), I7 =>  inp_feat(100)); 
C_30_S_3_L_5_inst : LUT8 generic map(INIT => "0011001011100010000000001000001101100000001100000000000000000010010000010000000000000000000100000000000000000000000000000000000010010010101100100010000000000000001110101010000000010100000000100000000000000010000100001000000000000000000000000000000000000000") port map( O =>C_30_S_3_L_5_out, I0 =>  inp_feat(468), I1 =>  inp_feat(394), I2 =>  inp_feat(477), I3 =>  inp_feat(275), I4 =>  inp_feat(508), I5 =>  inp_feat(120), I6 =>  inp_feat(393), I7 =>  inp_feat(344)); 
C_30_S_3_L_6_inst : LUT8 generic map(INIT => "1111000100110000101000001000000000000000101000000000000000000000111100001000000011000000100000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_3_L_6_out, I0 =>  inp_feat(469), I1 =>  inp_feat(509), I2 =>  inp_feat(100), I3 =>  inp_feat(262), I4 =>  inp_feat(58), I5 =>  inp_feat(64), I6 =>  inp_feat(18), I7 =>  inp_feat(341)); 
C_30_S_3_L_7_inst : LUT8 generic map(INIT => "1000100010000000010000000100000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000100011110100110000001100000011000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_3_L_7_out, I0 =>  inp_feat(120), I1 =>  inp_feat(477), I2 =>  inp_feat(474), I3 =>  inp_feat(124), I4 =>  inp_feat(458), I5 =>  inp_feat(258), I6 =>  inp_feat(393), I7 =>  inp_feat(277)); 
C_30_S_4_L_0_inst : LUT8 generic map(INIT => "0000001100000000100010000100010000001001000000001010110000000100001010000000000000000010010000000000000000000000000011101000100000000000000000000000100000000000000001000000000010001000010001000000000000000000110001000000000100000100000000001000010010001001") port map( O =>C_30_S_4_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(328), I2 =>  inp_feat(41), I3 =>  inp_feat(182), I4 =>  inp_feat(228), I5 =>  inp_feat(52), I6 =>  inp_feat(380), I7 =>  inp_feat(362)); 
C_30_S_4_L_1_inst : LUT8 generic map(INIT => "0000001000000010000000000000000010111000100000000000000000000000011000000110001010000000100010000000000010100000000000000000000011011010001000001000111011000000101100110011000000010000000000000000000000000000000000000000000000000000000000000000000000100000") port map( O =>C_30_S_4_L_1_out, I0 =>  inp_feat(353), I1 =>  inp_feat(120), I2 =>  inp_feat(420), I3 =>  inp_feat(82), I4 =>  inp_feat(413), I5 =>  inp_feat(144), I6 =>  inp_feat(74), I7 =>  inp_feat(95)); 
C_30_S_4_L_2_inst : LUT8 generic map(INIT => "1000001000001010000011110000000000000000000010000000000000000000000000100000000000001000000000000000000000000000000000000000000010101000000010001010101000000000101000000000000000000000100000001000001000100000000000000000000000000000000000000000000000000000") port map( O =>C_30_S_4_L_2_out, I0 =>  inp_feat(100), I1 =>  inp_feat(364), I2 =>  inp_feat(52), I3 =>  inp_feat(64), I4 =>  inp_feat(203), I5 =>  inp_feat(173), I6 =>  inp_feat(472), I7 =>  inp_feat(223)); 
C_30_S_4_L_3_inst : LUT8 generic map(INIT => "0000100000001000100000000000000000000000000000000000000000000000100110100100000100001010100111010000000000000000000000000000000011001000100010000000000000000000000010000000101000000000000000001000100010101010000000000000000010001000100010100000000000000000") port map( O =>C_30_S_4_L_3_out, I0 =>  inp_feat(449), I1 =>  inp_feat(261), I2 =>  inp_feat(29), I3 =>  inp_feat(119), I4 =>  inp_feat(331), I5 =>  inp_feat(8), I6 =>  inp_feat(56), I7 =>  inp_feat(223)); 
C_30_S_4_L_4_inst : LUT8 generic map(INIT => "1110011000000010010111010000000010010000000000101100100110001001010001001000001000000100100000001000101000000000000000000000100000000000000001000000110000000000000000000000000001000100000000001000010000000000000000000000100000000000000010100000000000000000") port map( O =>C_30_S_4_L_4_out, I0 =>  inp_feat(18), I1 =>  inp_feat(270), I2 =>  inp_feat(346), I3 =>  inp_feat(331), I4 =>  inp_feat(275), I5 =>  inp_feat(344), I6 =>  inp_feat(416), I7 =>  inp_feat(508)); 
C_30_S_4_L_5_inst : LUT8 generic map(INIT => "1111000000010000101100001010000001010000000000001011011000100000000000000000000001100100000000000000000000000000111100100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_30_S_4_L_5_out, I0 =>  inp_feat(283), I1 =>  inp_feat(291), I2 =>  inp_feat(57), I3 =>  inp_feat(506), I4 =>  inp_feat(61), I5 =>  inp_feat(256), I6 =>  inp_feat(174), I7 =>  inp_feat(393)); 
C_30_S_4_L_6_inst : LUT8 generic map(INIT => "0010100000000100100000000000100011000000000000000000000000000000001000000000001000000000000000000000000000100000000000000000000000101100000000000000101000000000101000000000000000000000000000001010100000001000001011000000100010000000000000000000000000100000") port map( O =>C_30_S_4_L_6_out, I0 =>  inp_feat(283), I1 =>  inp_feat(324), I2 =>  inp_feat(176), I3 =>  inp_feat(87), I4 =>  inp_feat(309), I5 =>  inp_feat(277), I6 =>  inp_feat(422), I7 =>  inp_feat(312)); 
C_30_S_4_L_7_inst : LUT8 generic map(INIT => "0011000001000000000000001000000000000000000000000000000000000000000100000111000000000000000000001000000010000000001000000000000011000010010011010011000001000000110000000100000000000000000000000100000011010000000000000100000011000000110000000000000000000000") port map( O =>C_30_S_4_L_7_out, I0 =>  inp_feat(460), I1 =>  inp_feat(198), I2 =>  inp_feat(351), I3 =>  inp_feat(291), I4 =>  inp_feat(326), I5 =>  inp_feat(124), I6 =>  inp_feat(434), I7 =>  inp_feat(178)); 
C_31_S_0_L_0_inst : LUT8 generic map(INIT => "1111101011111111100010001111000011010000110111111110101011110000110111101101000010000000000000000000000000110000100000000000000000000000000011011000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_31_S_0_L_0_out, I0 =>  inp_feat(141), I1 =>  inp_feat(201), I2 =>  inp_feat(459), I3 =>  inp_feat(472), I4 =>  inp_feat(167), I5 =>  inp_feat(221), I6 =>  inp_feat(157), I7 =>  inp_feat(299)); 
C_31_S_0_L_1_inst : LUT8 generic map(INIT => "0011111111000000111111001000000000101110100000001111000100000000110111111100000010000100000000001000000010000000000000000000000000100010110010000101110010001100001000011000110011001100000011001100111011001100110011001100110010001100110011000100110010001100") port map( O =>C_31_S_0_L_1_out, I0 =>  inp_feat(201), I1 =>  inp_feat(57), I2 =>  inp_feat(316), I3 =>  inp_feat(62), I4 =>  inp_feat(83), I5 =>  inp_feat(373), I6 =>  inp_feat(353), I7 =>  inp_feat(75)); 
C_31_S_0_L_2_inst : LUT8 generic map(INIT => "1001100011010000111100000000000010000000110000000100000000000000111011101000100011001100000000001100110000000000110001000000000011111000101000001101000000000000111100001110000000000000000000001010101010000000100000001000000010000000100000001000000010000000") port map( O =>C_31_S_0_L_2_out, I0 =>  inp_feat(304), I1 =>  inp_feat(223), I2 =>  inp_feat(29), I3 =>  inp_feat(238), I4 =>  inp_feat(37), I5 =>  inp_feat(256), I6 =>  inp_feat(98), I7 =>  inp_feat(197)); 
C_31_S_0_L_3_inst : LUT8 generic map(INIT => "1011000011100000111010101010111011000001010000001000000000000000101111101100100011101100110010001110110100000000101000000000000001001000110000101010000011100000111000101110000000000000000000001100100011001000111000001100010011101111000000000000000000000000") port map( O =>C_31_S_0_L_3_out, I0 =>  inp_feat(221), I1 =>  inp_feat(120), I2 =>  inp_feat(29), I3 =>  inp_feat(222), I4 =>  inp_feat(7), I5 =>  inp_feat(30), I6 =>  inp_feat(413), I7 =>  inp_feat(5)); 
C_31_S_0_L_4_inst : LUT8 generic map(INIT => "0011110111111101111111101100110100010000110011001011111011001100010011011100110000101101100001010000010101000000000011010000000100000000100000000100000000001100000000001000000001001000100000000000010100001100000011010000110000000001000000000000000000000000") port map( O =>C_31_S_0_L_4_out, I0 =>  inp_feat(71), I1 =>  inp_feat(111), I2 =>  inp_feat(187), I3 =>  inp_feat(336), I4 =>  inp_feat(316), I5 =>  inp_feat(31), I6 =>  inp_feat(115), I7 =>  inp_feat(144)); 
C_31_S_0_L_5_inst : LUT8 generic map(INIT => "0101110111101000110100110100000011101110111101000000101001100000000010001001100000000000100000000000000011110000100100000100000010101111100010001101100000000000100011001000000010000000000000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_31_S_0_L_5_out, I0 =>  inp_feat(206), I1 =>  inp_feat(373), I2 =>  inp_feat(98), I3 =>  inp_feat(459), I4 =>  inp_feat(221), I5 =>  inp_feat(176), I6 =>  inp_feat(464), I7 =>  inp_feat(366)); 
C_31_S_0_L_6_inst : LUT8 generic map(INIT => "0101000111011110010011011100100101000000110000001100000010000000110001001000010111000100110001000000000010000000110000001000000010000100110011001000110011001101000000000100000000000000000000000000000000000000000000000000010000000000000100000000000000000000") port map( O =>C_31_S_0_L_6_out, I0 =>  inp_feat(364), I1 =>  inp_feat(276), I2 =>  inp_feat(301), I3 =>  inp_feat(378), I4 =>  inp_feat(336), I5 =>  inp_feat(401), I6 =>  inp_feat(504), I7 =>  inp_feat(304)); 
C_31_S_0_L_7_inst : LUT8 generic map(INIT => "1110111110001111000000000000001010000101000011110000000000000000111010101000000010000010100000000000000010001000000000000000000000110011000010000000000000000000000000000000100000000000000000001100100010000000100000000000000000000000000000000000000000000000") port map( O =>C_31_S_0_L_7_out, I0 =>  inp_feat(211), I1 =>  inp_feat(249), I2 =>  inp_feat(419), I3 =>  inp_feat(501), I4 =>  inp_feat(300), I5 =>  inp_feat(18), I6 =>  inp_feat(306), I7 =>  inp_feat(256)); 
C_31_S_1_L_0_inst : LUT8 generic map(INIT => "1111110011011100111000001000000011111100110111001110100011011000010111000101010111101100010101001100010001011100010001000000010001010000110101000111000010000000011101001101000001110000111100000101000001010100111101000101000000100000010000001111110001010100") port map( O =>C_31_S_1_L_0_out, I0 =>  inp_feat(239), I1 =>  inp_feat(178), I2 =>  inp_feat(222), I3 =>  inp_feat(193), I4 =>  inp_feat(413), I5 =>  inp_feat(362), I6 =>  inp_feat(52), I7 =>  inp_feat(29)); 
C_31_S_1_L_1_inst : LUT8 generic map(INIT => "0111110111101010001101001000000001111111101010100000010010000000101000100010101010110101000000001110111010101010000000000000000001000000110010100000000000000000001000001000101000000000000000000000001000101010000000000000000010001010101010100000000000000000") port map( O =>C_31_S_1_L_1_out, I0 =>  inp_feat(30), I1 =>  inp_feat(336), I2 =>  inp_feat(283), I3 =>  inp_feat(98), I4 =>  inp_feat(339), I5 =>  inp_feat(328), I6 =>  inp_feat(304), I7 =>  inp_feat(460)); 
C_31_S_1_L_2_inst : LUT8 generic map(INIT => "1111110100000100001111111110010111111111101010001111111110101111011010001000100011111111111011101100000010000000111111110111111100000000100000000010000110011110001001010010100000100101001110111000001110101000111111111111111010000000100000001111111111111111") port map( O =>C_31_S_1_L_2_out, I0 =>  inp_feat(83), I1 =>  inp_feat(201), I2 =>  inp_feat(41), I3 =>  inp_feat(451), I4 =>  inp_feat(182), I5 =>  inp_feat(420), I6 =>  inp_feat(82), I7 =>  inp_feat(221)); 
C_31_S_1_L_3_inst : LUT8 generic map(INIT => "0000010011111101000001010111110101000100110100000000000011001001111011001100110111101101110001000100000001001100000000000000010011001100110111011101110111010100000000001100010000000000000011011100110011011100011001010101010100000000000011000000000000000100") port map( O =>C_31_S_1_L_3_out, I0 =>  inp_feat(141), I1 =>  inp_feat(339), I2 =>  inp_feat(259), I3 =>  inp_feat(62), I4 =>  inp_feat(373), I5 =>  inp_feat(144), I6 =>  inp_feat(161), I7 =>  inp_feat(498)); 
C_31_S_1_L_4_inst : LUT8 generic map(INIT => "1011111011110100000011010000010010000000001000101000100000000000100011000000000010101000000000001010111000100010101011000000000000011000001111000000000000000101000000110000000000000000000000001010111100000000000000000000000000100010000000000000000100000000") port map( O =>C_31_S_1_L_4_out, I0 =>  inp_feat(46), I1 =>  inp_feat(71), I2 =>  inp_feat(364), I3 =>  inp_feat(74), I4 =>  inp_feat(233), I5 =>  inp_feat(256), I6 =>  inp_feat(264), I7 =>  inp_feat(52)); 
C_31_S_1_L_5_inst : LUT8 generic map(INIT => "0100101011010111010110101111000011011010100010000000000000000000010010000000000000100000000000001110101000000000001000100000000001001100110011110000000011000000011100101100101000110000010000000000000000001000100000000000000000000000000000000010000000000000") port map( O =>C_31_S_1_L_5_out, I0 =>  inp_feat(331), I1 =>  inp_feat(328), I2 =>  inp_feat(84), I3 =>  inp_feat(354), I4 =>  inp_feat(15), I5 =>  inp_feat(419), I6 =>  inp_feat(229), I7 =>  inp_feat(82)); 
C_31_S_1_L_6_inst : LUT8 generic map(INIT => "1111100111101110110111100010000001110101110000001000100010101010000100001100010000000000000000000100000000000000000000000010000011110101110000011110000000100000001000001000000010100010101010100101010001000000001000000000000000000000000000000010001010100010") port map( O =>C_31_S_1_L_6_out, I0 =>  inp_feat(200), I1 =>  inp_feat(504), I2 =>  inp_feat(31), I3 =>  inp_feat(344), I4 =>  inp_feat(332), I5 =>  inp_feat(229), I6 =>  inp_feat(5), I7 =>  inp_feat(141)); 
C_31_S_1_L_7_inst : LUT8 generic map(INIT => "0000110011111111100010000000110001101000111110101010000000101000000011001110101010001000000010001010001000001111100011000000111111000000111111110000000010001111110000001111111110000000101011110000000001000110000000001000111000000000001011110000000010001111") port map( O =>C_31_S_1_L_7_out, I0 =>  inp_feat(339), I1 =>  inp_feat(52), I2 =>  inp_feat(390), I3 =>  inp_feat(354), I4 =>  inp_feat(259), I5 =>  inp_feat(420), I6 =>  inp_feat(373), I7 =>  inp_feat(353)); 
C_31_S_2_L_0_inst : LUT8 generic map(INIT => "1111111111101010000011011100000011101110110000100000000000000000011000101110000000000000110000001110000010000000000000000000000010001000101010100000000100000000000000000000000000000010000000000000001010101010000000000000000000000000101100100000000000000000") port map( O =>C_31_S_2_L_0_out, I0 =>  inp_feat(5), I1 =>  inp_feat(51), I2 =>  inp_feat(139), I3 =>  inp_feat(98), I4 =>  inp_feat(464), I5 =>  inp_feat(256), I6 =>  inp_feat(157), I7 =>  inp_feat(29)); 
C_31_S_2_L_1_inst : LUT8 generic map(INIT => "1111111100000000111111000000000011111100100000001111110001010100110000000000000001010100000000001101000000000000011000000000000000011001000000001100000000000000101010000000100000000000000000000101100000000000010001000000000000000000000000000000000000000000") port map( O =>C_31_S_2_L_1_out, I0 =>  inp_feat(248), I1 =>  inp_feat(41), I2 =>  inp_feat(428), I3 =>  inp_feat(18), I4 =>  inp_feat(82), I5 =>  inp_feat(316), I6 =>  inp_feat(339), I7 =>  inp_feat(256)); 
C_31_S_2_L_2_inst : LUT8 generic map(INIT => "1111000011110000001000000010000010000000011000001010000010100000111010001111000000100000111100001010000011110010101000101111000000100000101100001000001010100000001000001010000000100000100000000100000011110000001000101111000000100000001100001010000011111000") port map( O =>C_31_S_2_L_2_out, I0 =>  inp_feat(144), I1 =>  inp_feat(316), I2 =>  inp_feat(299), I3 =>  inp_feat(182), I4 =>  inp_feat(161), I5 =>  inp_feat(373), I6 =>  inp_feat(362), I7 =>  inp_feat(52)); 
C_31_S_2_L_3_inst : LUT8 generic map(INIT => "0100100000000000111101001100010100000100000010001111010101000101010110000000000001010100010100001100000001010000010101000101010001011000000000001101010101010100110000001000000001010100010001001100100010100000010101011101010001000000011101000101010101010101") port map( O =>C_31_S_2_L_3_out, I0 =>  inp_feat(413), I1 =>  inp_feat(29), I2 =>  inp_feat(196), I3 =>  inp_feat(174), I4 =>  inp_feat(98), I5 =>  inp_feat(265), I6 =>  inp_feat(304), I7 =>  inp_feat(328)); 
C_31_S_2_L_4_inst : LUT8 generic map(INIT => "0010101111111011100010011101110100001000000000000000110011001100101111110000100011001101000000000000100000000000000010000000000010101000101010000000100010001000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_31_S_2_L_4_out, I0 =>  inp_feat(229), I1 =>  inp_feat(98), I2 =>  inp_feat(4), I3 =>  inp_feat(328), I4 =>  inp_feat(419), I5 =>  inp_feat(249), I6 =>  inp_feat(206), I7 =>  inp_feat(20)); 
C_31_S_2_L_5_inst : LUT8 generic map(INIT => "1111101101100010001100101111000011110111111100001111001010110000111100111001000000100000110000001111010111110000011100001111000011000000100100001000001001110000111100000011000000010000001100001111001011100000101000100110000001010000111100000001000011110000") port map( O =>C_31_S_2_L_5_out, I0 =>  inp_feat(500), I1 =>  inp_feat(362), I2 =>  inp_feat(97), I3 =>  inp_feat(210), I4 =>  inp_feat(373), I5 =>  inp_feat(353), I6 =>  inp_feat(52), I7 =>  inp_feat(161)); 
C_31_S_2_L_6_inst : LUT8 generic map(INIT => "0111001010101000110100000101000001110000111100100011000011100000111000000111000000000000110100000000000010000000000000001000000011100000110000001010000010010000000000001000000010001000100000000000000010000000101000001111000000000000000000000000000000000000") port map( O =>C_31_S_2_L_6_out, I0 =>  inp_feat(480), I1 =>  inp_feat(290), I2 =>  inp_feat(299), I3 =>  inp_feat(161), I4 =>  inp_feat(83), I5 =>  inp_feat(485), I6 =>  inp_feat(492), I7 =>  inp_feat(186)); 
C_31_S_2_L_7_inst : LUT8 generic map(INIT => "1100000111110000110000001000000011010001111110000000000010001000111100011001001100000000000000001100001011111010000000001010000011100100110100000000000010000000010100001010100000000000000000000000000010100000000000000000000000100010111110100000000000000000") port map( O =>C_31_S_2_L_7_out, I0 =>  inp_feat(198), I1 =>  inp_feat(229), I2 =>  inp_feat(460), I3 =>  inp_feat(413), I4 =>  inp_feat(144), I5 =>  inp_feat(346), I6 =>  inp_feat(102), I7 =>  inp_feat(52)); 
C_31_S_3_L_0_inst : LUT8 generic map(INIT => "0100000011000000111011100000000011000000010000001100110000000000110010001000000000000000000000001000000000000000000000000000000011111010100000001000101000000000101010000000000000000000000000001010100000000000000000000000000010001000000000000000000000000000") port map( O =>C_31_S_3_L_0_out, I0 =>  inp_feat(475), I1 =>  inp_feat(37), I2 =>  inp_feat(491), I3 =>  inp_feat(339), I4 =>  inp_feat(395), I5 =>  inp_feat(337), I6 =>  inp_feat(238), I7 =>  inp_feat(306)); 
C_31_S_3_L_1_inst : LUT8 generic map(INIT => "1111110011110000111010000000000000100000100000001000100000000000101110100100000011001100000010000101100000000000000000000000000011001100000000001100110000000000000000000000000000000000000000000111110101100000110011000000000000000000000000000000000000000000") port map( O =>C_31_S_3_L_1_out, I0 =>  inp_feat(378), I1 =>  inp_feat(75), I2 =>  inp_feat(265), I3 =>  inp_feat(500), I4 =>  inp_feat(308), I5 =>  inp_feat(360), I6 =>  inp_feat(221), I7 =>  inp_feat(304)); 
C_31_S_3_L_2_inst : LUT8 generic map(INIT => "0010111001001100110010001100100000001000000010000000100000001000000010001100100010001000100000000000000000000000000000000000000011011100010111001000100000001000101110101100101000001000000010001000000011011100100010001100100010101010000010100000000000000000") port map( O =>C_31_S_3_L_2_out, I0 =>  inp_feat(323), I1 =>  inp_feat(300), I2 =>  inp_feat(295), I3 =>  inp_feat(303), I4 =>  inp_feat(470), I5 =>  inp_feat(144), I6 =>  inp_feat(52), I7 =>  inp_feat(141)); 
C_31_S_3_L_3_inst : LUT8 generic map(INIT => "1010111011101111101011100000001110001010111110111000101010111111011000001101011000000000011000000000000001010001000000001000000111100000111100000010100010110011100000001111000010101000101100111111000011110101110000000110001100100000101100010000000000110011") port map( O =>C_31_S_3_L_3_out, I0 =>  inp_feat(221), I1 =>  inp_feat(81), I2 =>  inp_feat(378), I3 =>  inp_feat(357), I4 =>  inp_feat(37), I5 =>  inp_feat(322), I6 =>  inp_feat(256), I7 =>  inp_feat(87)); 
C_31_S_3_L_4_inst : LUT8 generic map(INIT => "0010111111101011110011011111010110000000111000010000000011110101100011110000000110000101000001011001000000000001000001010000010100001001111010000000000101010100000000000000010000000000000101011100110101010101100001010000010100000101000001010000010100000101") port map( O =>C_31_S_3_L_4_out, I0 =>  inp_feat(346), I1 =>  inp_feat(37), I2 =>  inp_feat(232), I3 =>  inp_feat(143), I4 =>  inp_feat(187), I5 =>  inp_feat(304), I6 =>  inp_feat(87), I7 =>  inp_feat(229)); 
C_31_S_3_L_5_inst : LUT8 generic map(INIT => "0111111110111111010101110011000100110010001010111011001001000000100000011101011001011111010001100100000000010111100101000000000001011111110111111101111011010111110101010101010001110100010100000100000001000111110111111101110101001100010101001100100001000100") port map( O =>C_31_S_3_L_5_out, I0 =>  inp_feat(336), I1 =>  inp_feat(331), I2 =>  inp_feat(316), I3 =>  inp_feat(500), I4 =>  inp_feat(451), I5 =>  inp_feat(339), I6 =>  inp_feat(41), I7 =>  inp_feat(82)); 
C_31_S_3_L_6_inst : LUT8 generic map(INIT => "0101110111111011011100111100101010100000110010000001101011001110101010100011001000000101111000100000000010001100000000001000000000001000100011101111011111110110100000001100101011011001110011111000110011000110011000100110111110001000110010001100000011001100") port map( O =>C_31_S_3_L_6_out, I0 =>  inp_feat(451), I1 =>  inp_feat(220), I2 =>  inp_feat(373), I3 =>  inp_feat(336), I4 =>  inp_feat(210), I5 =>  inp_feat(148), I6 =>  inp_feat(120), I7 =>  inp_feat(141)); 
C_31_S_3_L_7_inst : LUT8 generic map(INIT => "1111111101010010001001110011000100001010111100000000001000000000111100101111001001110010001000111000001001110000000000000000000000100011000000110000001100001011000000000011100000000000000000100000001100010000000000110001001100000000000000000000001000000000") port map( O =>C_31_S_3_L_7_out, I0 =>  inp_feat(301), I1 =>  inp_feat(4), I2 =>  inp_feat(351), I3 =>  inp_feat(373), I4 =>  inp_feat(238), I5 =>  inp_feat(342), I6 =>  inp_feat(290), I7 =>  inp_feat(256)); 
C_31_S_4_L_0_inst : LUT8 generic map(INIT => "1101111111110110111101111000001001110011000000001111111010100000111110100011000010110010001100100000000000000000101000000000000001000010000001001101110011010100010000000000000011010100000000000000010100000100100000100100010000000000000000000000000100000001") port map( O =>C_31_S_4_L_0_out, I0 =>  inp_feat(61), I1 =>  inp_feat(329), I2 =>  inp_feat(201), I3 =>  inp_feat(228), I4 =>  inp_feat(336), I5 =>  inp_feat(130), I6 =>  inp_feat(71), I7 =>  inp_feat(157)); 
C_31_S_4_L_1_inst : LUT8 generic map(INIT => "0111111000011110011000101000000011101010111110101000000001000000001000101000101000100010000000101000100010001000000000001000100010101000100010000000000010000000101010001000100000001000100010000000000010000000000000000000000010101000100010001000000010000000") port map( O =>C_31_S_4_L_1_out, I0 =>  inp_feat(30), I1 =>  inp_feat(354), I2 =>  inp_feat(378), I3 =>  inp_feat(468), I4 =>  inp_feat(256), I5 =>  inp_feat(98), I6 =>  inp_feat(157), I7 =>  inp_feat(309)); 
C_31_S_4_L_2_inst : LUT8 generic map(INIT => "1101110001001100111100000001000001111100001000001011000000110000010111100110011001111110000110101011000000110000111101000011000011000100010101001000000000000000100000000000000010000000001100000000010010101100001000000000000000000000001100000000000000100000") port map( O =>C_31_S_4_L_2_out, I0 =>  inp_feat(331), I1 =>  inp_feat(302), I2 =>  inp_feat(346), I3 =>  inp_feat(29), I4 =>  inp_feat(290), I5 =>  inp_feat(374), I6 =>  inp_feat(413), I7 =>  inp_feat(470)); 
C_31_S_4_L_3_inst : LUT8 generic map(INIT => "1010111110101000001001000000100001110111011100001011110010110000000001010000111100100111001111110011111101000100000111110011001111001000100010000000000010001000010101000000000000000100000000000001011111111000010101110011000100110111011100000111011100110001") port map( O =>C_31_S_4_L_3_out, I0 =>  inp_feat(307), I1 =>  inp_feat(336), I2 =>  inp_feat(328), I3 =>  inp_feat(378), I4 =>  inp_feat(304), I5 =>  inp_feat(265), I6 =>  inp_feat(52), I7 =>  inp_feat(342)); 
C_31_S_4_L_4_inst : LUT8 generic map(INIT => "1011101010001101111111010001100101000001000000001100110000000000110011000000010010000000000000000000000000000000000000000000000000000000000001001000101000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_31_S_4_L_4_out, I0 =>  inp_feat(201), I1 =>  inp_feat(339), I2 =>  inp_feat(58), I3 =>  inp_feat(95), I4 =>  inp_feat(336), I5 =>  inp_feat(464), I6 =>  inp_feat(342), I7 =>  inp_feat(299)); 
C_31_S_4_L_5_inst : LUT8 generic map(INIT => "1101110001101011001101110000110011111010000000110010110100000010010011100000001011001111100001011100011000000000100010110000110011110000001000001001101010011010101000000010001000000000100000101100100010000000110011111000111111001000110010001000100010001011") port map( O =>C_31_S_4_L_5_out, I0 =>  inp_feat(109), I1 =>  inp_feat(220), I2 =>  inp_feat(53), I3 =>  inp_feat(52), I4 =>  inp_feat(210), I5 =>  inp_feat(120), I6 =>  inp_feat(141), I7 =>  inp_feat(353)); 
C_31_S_4_L_6_inst : LUT8 generic map(INIT => "1011101011101000101010001110000011111011101110110111101110111011111110001010100000101000101000001001000010001000101010000010100000100010010010000000100000001000001000100000100000110010001110100000000000001000000000000000000000110000000010000000000010001000") port map( O =>C_31_S_4_L_6_out, I0 =>  inp_feat(256), I1 =>  inp_feat(98), I2 =>  inp_feat(328), I3 =>  inp_feat(378), I4 =>  inp_feat(3), I5 =>  inp_feat(273), I6 =>  inp_feat(198), I7 =>  inp_feat(211)); 
C_31_S_4_L_7_inst : LUT8 generic map(INIT => "0111001000100010101100001010000011100010010000100000000010000000101000100010100010100000000000100000001000000000000000000000000011111111101111111010000000000010100010001110001010000000100000000011101100111001111100000001000010000010000000110000000010000000") port map( O =>C_31_S_4_L_7_out, I0 =>  inp_feat(306), I1 =>  inp_feat(98), I2 =>  inp_feat(274), I3 =>  inp_feat(29), I4 =>  inp_feat(198), I5 =>  inp_feat(302), I6 =>  inp_feat(229), I7 =>  inp_feat(413)); 
C_32_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_0_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_1_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_2_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_3_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_4_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_5_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_6_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_0_L_7_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_0_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_1_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_2_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_3_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_4_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_5_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_6_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_1_L_7_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_0_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_1_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_2_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_3_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_4_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_5_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_6_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_2_L_7_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_0_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_1_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_2_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_3_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_4_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_5_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_6_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_3_L_7_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_0_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_1_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_2_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_3_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_4_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_5_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_6_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_32_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000001000000010001000100010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000001010101010100000") port map( O =>C_32_S_4_L_7_out, I0 =>  inp_feat(9), I1 =>  inp_feat(222), I2 =>  inp_feat(179), I3 =>  inp_feat(466), I4 =>  inp_feat(161), I5 =>  inp_feat(48), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_33_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000010000000100000000000000000000000000000000000000000000000000000000001011010111000010110000000000000000100100000000000000000000000000000101000000000000000000000000000000000000000000000001000000000000010101010000000000000000000000000000000000000000") port map( O =>C_33_S_0_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(310), I2 =>  inp_feat(367), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_33_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000001000000100000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000010110000001100010011110111111000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_0_L_1_out, I0 =>  inp_feat(298), I1 =>  inp_feat(367), I2 =>  inp_feat(382), I3 =>  inp_feat(469), I4 =>  inp_feat(218), I5 =>  inp_feat(286), I6 =>  inp_feat(26), I7 =>  inp_feat(509)); 
C_33_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000001000000000000011100000000000010000000010000010101000000000000001000000000000000110000000000000100000000000100001000000001000001010000000100000101000000000100110100000000010001010001000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_0_L_2_out, I0 =>  inp_feat(382), I1 =>  inp_feat(7), I2 =>  inp_feat(48), I3 =>  inp_feat(509), I4 =>  inp_feat(273), I5 =>  inp_feat(301), I6 =>  inp_feat(147), I7 =>  inp_feat(373)); 
C_33_S_0_L_3_inst : LUT8 generic map(INIT => "0000000001000000000000000000000100000000000000100000101000010011000000000000000000000000000000000000000000000000000000000000000001000001000111110000101110110111000000000000111100000000000111110000000000000000000100010001000000000000000000000000000000000000") port map( O =>C_33_S_0_L_3_out, I0 =>  inp_feat(469), I1 =>  inp_feat(218), I2 =>  inp_feat(435), I3 =>  inp_feat(303), I4 =>  inp_feat(494), I5 =>  inp_feat(244), I6 =>  inp_feat(213), I7 =>  inp_feat(310)); 
C_33_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011000000010010001100000001010001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_0_L_4_out, I0 =>  inp_feat(420), I1 =>  inp_feat(416), I2 =>  inp_feat(178), I3 =>  inp_feat(19), I4 =>  inp_feat(364), I5 =>  inp_feat(237), I6 =>  inp_feat(26), I7 =>  inp_feat(218)); 
C_33_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010001001000000100000000000000000011000110000000000000000000000001111111101100010000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001110001000000000000000000000000") port map( O =>C_33_S_0_L_5_out, I0 =>  inp_feat(7), I1 =>  inp_feat(303), I2 =>  inp_feat(247), I3 =>  inp_feat(9), I4 =>  inp_feat(495), I5 =>  inp_feat(142), I6 =>  inp_feat(218), I7 =>  inp_feat(466)); 
C_33_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000001101000000000000000010111011000010110000000000000000000000000000000000000010000000000000001100001001000000000000000010000000000001010000000000000000001010100000111100000000000000000000000000000000000000000000000000100011000000110000000000000000") port map( O =>C_33_S_0_L_6_out, I0 =>  inp_feat(373), I1 =>  inp_feat(469), I2 =>  inp_feat(382), I3 =>  inp_feat(247), I4 =>  inp_feat(26), I5 =>  inp_feat(218), I6 =>  inp_feat(362), I7 =>  inp_feat(57)); 
C_33_S_0_L_7_inst : LUT8 generic map(INIT => "0000001000000100000000000000000000000010000000101010101000000010000000000000000000000000000000000000000000000000000000000000000000100001000000001010001000000000000000000000000110101010101010100000000000000010000000000000000000000000000000000000000010001100") port map( O =>C_33_S_0_L_7_out, I0 =>  inp_feat(180), I1 =>  inp_feat(53), I2 =>  inp_feat(469), I3 =>  inp_feat(356), I4 =>  inp_feat(48), I5 =>  inp_feat(77), I6 =>  inp_feat(464), I7 =>  inp_feat(212)); 
C_33_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000010000000100000000000000000000000000000000000000000000000000000000001011010111000010110000000000000000100100000000000000000000000000000101000000000000000000000000000000000000000000000001000000000000010101010000000000000000000000000000000000000000") port map( O =>C_33_S_1_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(310), I2 =>  inp_feat(367), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_33_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000001000000100000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000010110000001100010011110111111000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_1_L_1_out, I0 =>  inp_feat(298), I1 =>  inp_feat(367), I2 =>  inp_feat(382), I3 =>  inp_feat(469), I4 =>  inp_feat(218), I5 =>  inp_feat(286), I6 =>  inp_feat(26), I7 =>  inp_feat(509)); 
C_33_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000001000000101100000000000000000000001100000000000000000000110000000000000011000000000000010000000000100000000100000000000010000000010000001100000000000000000000000000100000000000100001001001000000000000110000000000010000000000000000000000") port map( O =>C_33_S_1_L_2_out, I0 =>  inp_feat(88), I1 =>  inp_feat(112), I2 =>  inp_feat(48), I3 =>  inp_feat(142), I4 =>  inp_feat(386), I5 =>  inp_feat(200), I6 =>  inp_feat(301), I7 =>  inp_feat(19)); 
C_33_S_1_L_3_inst : LUT8 generic map(INIT => "0001000000101100000000000000000000000101011001010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_1_L_3_out, I0 =>  inp_feat(382), I1 =>  inp_feat(256), I2 =>  inp_feat(420), I3 =>  inp_feat(52), I4 =>  inp_feat(119), I5 =>  inp_feat(303), I6 =>  inp_feat(26), I7 =>  inp_feat(9)); 
C_33_S_1_L_4_inst : LUT8 generic map(INIT => "0000010000000000010001010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000011001100100010000100110000000000000000000000000011000000000000000000100000001000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_1_L_4_out, I0 =>  inp_feat(157), I1 =>  inp_feat(178), I2 =>  inp_feat(303), I3 =>  inp_feat(154), I4 =>  inp_feat(242), I5 =>  inp_feat(216), I6 =>  inp_feat(92), I7 =>  inp_feat(161)); 
C_33_S_1_L_5_inst : LUT8 generic map(INIT => "0000001000000000000100000000000000010011000000000011000100000000000100000000000000010010000100000101001100000000000100010001000000000000000000000000000000000000000000000000000001010000000000000100000000000000000000000000000000010001000000000001000100010000") port map( O =>C_33_S_1_L_5_out, I0 =>  inp_feat(382), I1 =>  inp_feat(509), I2 =>  inp_feat(136), I3 =>  inp_feat(154), I4 =>  inp_feat(301), I5 =>  inp_feat(218), I6 =>  inp_feat(310), I7 =>  inp_feat(370)); 
C_33_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000010000000000000010000000000001000000000000000000000000000000100000000000100100000000000000000000000000001000110011000000000011001100000011001100010001000000110000000000000000000000000000000000000000001010100000001100000001000000") port map( O =>C_33_S_1_L_6_out, I0 =>  inp_feat(212), I1 =>  inp_feat(389), I2 =>  inp_feat(98), I3 =>  inp_feat(19), I4 =>  inp_feat(406), I5 =>  inp_feat(367), I6 =>  inp_feat(156), I7 =>  inp_feat(218)); 
C_33_S_1_L_7_inst : LUT8 generic map(INIT => "0011000000100000001000110000001001010101000000000100010100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001111100000000000000010000000000000111000000000000000000000000000000000000000000000000000000000000001000000000") port map( O =>C_33_S_1_L_7_out, I0 =>  inp_feat(48), I1 =>  inp_feat(310), I2 =>  inp_feat(303), I3 =>  inp_feat(215), I4 =>  inp_feat(247), I5 =>  inp_feat(207), I6 =>  inp_feat(286), I7 =>  inp_feat(480)); 
C_33_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000010000000100000000000000000000000000000000000000000000000000000000001011010111000010110000000000000000100100000000000000000000000000000101000000000000000000000000000000000000000000000001000000000000010101010000000000000000000000000000000000000000") port map( O =>C_33_S_2_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(310), I2 =>  inp_feat(367), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_33_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000001000000100000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000010110000001100010011110111111000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_2_L_1_out, I0 =>  inp_feat(298), I1 =>  inp_feat(367), I2 =>  inp_feat(382), I3 =>  inp_feat(469), I4 =>  inp_feat(218), I5 =>  inp_feat(286), I6 =>  inp_feat(26), I7 =>  inp_feat(509)); 
C_33_S_2_L_2_inst : LUT8 generic map(INIT => "0000000100000000000100010000000000000010000000000000000100000000000100000000000000010001000000000000000000000000000000110000000000000000000100000011000000000000000010000000000000000000000000000101000000000001011100010000000000000000010000001100000000000000") port map( O =>C_33_S_2_L_2_out, I0 =>  inp_feat(218), I1 =>  inp_feat(48), I2 =>  inp_feat(455), I3 =>  inp_feat(178), I4 =>  inp_feat(161), I5 =>  inp_feat(200), I6 =>  inp_feat(301), I7 =>  inp_feat(19)); 
C_33_S_2_L_3_inst : LUT8 generic map(INIT => "0000110001101111000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_2_L_3_out, I0 =>  inp_feat(257), I1 =>  inp_feat(373), I2 =>  inp_feat(420), I3 =>  inp_feat(303), I4 =>  inp_feat(83), I5 =>  inp_feat(26), I6 =>  inp_feat(234), I7 =>  inp_feat(444)); 
C_33_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010110000011101110000000000110000010000000000000011000000000000000000000000000000000000000000000001000000000000000000000000000000") port map( O =>C_33_S_2_L_4_out, I0 =>  inp_feat(86), I1 =>  inp_feat(19), I2 =>  inp_feat(115), I3 =>  inp_feat(364), I4 =>  inp_feat(117), I5 =>  inp_feat(425), I6 =>  inp_feat(216), I7 =>  inp_feat(218)); 
C_33_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000100000000000001000000000000000001000000000000000000000000010001010000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000101010101010000000001010101000000000000000000000000010001000") port map( O =>C_33_S_2_L_5_out, I0 =>  inp_feat(103), I1 =>  inp_feat(466), I2 =>  inp_feat(127), I3 =>  inp_feat(509), I4 =>  inp_feat(186), I5 =>  inp_feat(347), I6 =>  inp_feat(161), I7 =>  inp_feat(257)); 
C_33_S_2_L_6_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000000000000011000000000010000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000100100010001100110001000000010001000100000000000000000000000000100000000000010000000100000001000100") port map( O =>C_33_S_2_L_6_out, I0 =>  inp_feat(298), I1 =>  inp_feat(314), I2 =>  inp_feat(367), I3 =>  inp_feat(77), I4 =>  inp_feat(37), I5 =>  inp_feat(161), I6 =>  inp_feat(254), I7 =>  inp_feat(142)); 
C_33_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000010100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100100110000001001110011000000000000000000000011000000010000000000000000000000000000001100000000000000000000000000000000") port map( O =>C_33_S_2_L_7_out, I0 =>  inp_feat(303), I1 =>  inp_feat(509), I2 =>  inp_feat(494), I3 =>  inp_feat(382), I4 =>  inp_feat(218), I5 =>  inp_feat(17), I6 =>  inp_feat(20), I7 =>  inp_feat(142)); 
C_33_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000010000000100000000000000000000000000000000000000000000000000000000001011010111000010110000000000000000100100000000000000000000000000000101000000000000000000000000000000000000000000000001000000000000010101010000000000000000000000000000000000000000") port map( O =>C_33_S_3_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(310), I2 =>  inp_feat(367), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_33_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001001000000000000000000000000000001000000000000000000000000000000000000000000000000000011000001101101010100000000101000000000100011111111000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_3_L_1_out, I0 =>  inp_feat(310), I1 =>  inp_feat(333), I2 =>  inp_feat(227), I3 =>  inp_feat(151), I4 =>  inp_feat(382), I5 =>  inp_feat(121), I6 =>  inp_feat(26), I7 =>  inp_feat(509)); 
C_33_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000001010100000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010101010001000101010101010101010000000000000000000000000101111100000000000000000000000000010000000000000000000000000000000100000") port map( O =>C_33_S_3_L_2_out, I0 =>  inp_feat(390), I1 =>  inp_feat(469), I2 =>  inp_feat(247), I3 =>  inp_feat(88), I4 =>  inp_feat(310), I5 =>  inp_feat(154), I6 =>  inp_feat(286), I7 =>  inp_feat(52)); 
C_33_S_3_L_3_inst : LUT8 generic map(INIT => "0000000100011001000000000011000100000100100000000000000000000000000000000000000000000000000000000000000000001000000010000000000000100000001000110111000000110011000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000") port map( O =>C_33_S_3_L_3_out, I0 =>  inp_feat(434), I1 =>  inp_feat(382), I2 =>  inp_feat(86), I3 =>  inp_feat(161), I4 =>  inp_feat(212), I5 =>  inp_feat(271), I6 =>  inp_feat(331), I7 =>  inp_feat(301)); 
C_33_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000111000000000000000000000001000000010000000000000000000000111000010100000000000000000000000000000000000000000000110010000100000011110000000000000000000000100000000100000000000010000000101100001011000000000000000000000000000000000000") port map( O =>C_33_S_3_L_4_out, I0 =>  inp_feat(301), I1 =>  inp_feat(170), I2 =>  inp_feat(286), I3 =>  inp_feat(247), I4 =>  inp_feat(509), I5 =>  inp_feat(464), I6 =>  inp_feat(136), I7 =>  inp_feat(207)); 
C_33_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000010000000100000000000000010000000000000000000000000000000000000100000001010000000000000101000000011000000001000000000000000000011100000101100000000000010100000") port map( O =>C_33_S_3_L_5_out, I0 =>  inp_feat(286), I1 =>  inp_feat(373), I2 =>  inp_feat(26), I3 =>  inp_feat(142), I4 =>  inp_feat(396), I5 =>  inp_feat(509), I6 =>  inp_feat(469), I7 =>  inp_feat(310)); 
C_33_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010001000010000000000010011100101110001000000000001000101011111000100110010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000001000000001000100") port map( O =>C_33_S_3_L_6_out, I0 =>  inp_feat(247), I1 =>  inp_feat(56), I2 =>  inp_feat(186), I3 =>  inp_feat(406), I4 =>  inp_feat(218), I5 =>  inp_feat(469), I6 =>  inp_feat(382), I7 =>  inp_feat(474)); 
C_33_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000010000000000000000000001000001000000000000000000000000100100101001100001000000000100000001011110011001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000100000000000") port map( O =>C_33_S_3_L_7_out, I0 =>  inp_feat(470), I1 =>  inp_feat(161), I2 =>  inp_feat(86), I3 =>  inp_feat(303), I4 =>  inp_feat(466), I5 =>  inp_feat(469), I6 =>  inp_feat(509), I7 =>  inp_feat(12)); 
C_33_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000010000000100000000000000000000000000000000000000000000000000000000001011010111000010110000000000000000100100000000000000000000000000000101000000000000000000000000000000000000000000000001000000000000010101010000000000000000000000000000000000000000") port map( O =>C_33_S_4_L_0_out, I0 =>  inp_feat(382), I1 =>  inp_feat(310), I2 =>  inp_feat(367), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_33_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001001000000000000000000000000000001000000000000000000000000000000000000000000000000000011000001101101010100000000101000000000100011111111000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_4_L_1_out, I0 =>  inp_feat(310), I1 =>  inp_feat(333), I2 =>  inp_feat(227), I3 =>  inp_feat(151), I4 =>  inp_feat(382), I5 =>  inp_feat(121), I6 =>  inp_feat(26), I7 =>  inp_feat(509)); 
C_33_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000001010100000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010101010001000101010101010101010000000000000000000000000101111100000000000000000000000000010000000000000000000000000000000100000") port map( O =>C_33_S_4_L_2_out, I0 =>  inp_feat(390), I1 =>  inp_feat(469), I2 =>  inp_feat(247), I3 =>  inp_feat(88), I4 =>  inp_feat(310), I5 =>  inp_feat(154), I6 =>  inp_feat(286), I7 =>  inp_feat(52)); 
C_33_S_4_L_3_inst : LUT8 generic map(INIT => "0000001010010000001000000011000000000000110000000000000000000000000000000000000000000000000100000000000010000000000000000000000010110000001100001011000000110000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000") port map( O =>C_33_S_4_L_3_out, I0 =>  inp_feat(88), I1 =>  inp_feat(382), I2 =>  inp_feat(26), I3 =>  inp_feat(333), I4 =>  inp_feat(303), I5 =>  inp_feat(271), I6 =>  inp_feat(331), I7 =>  inp_feat(301)); 
C_33_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000001110010000000000000001000000000000000000000000000000000000000000000000000000000001000000000000011110000000000000000000000000000111100000000000000010000000000000000000000000000000000000000000001010000000000000000000000000000") port map( O =>C_33_S_4_L_4_out, I0 =>  inp_feat(386), I1 =>  inp_feat(302), I2 =>  inp_feat(111), I3 =>  inp_feat(119), I4 =>  inp_feat(180), I5 =>  inp_feat(19), I6 =>  inp_feat(12), I7 =>  inp_feat(86)); 
C_33_S_4_L_5_inst : LUT8 generic map(INIT => "0000001000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011101011110000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_4_L_5_out, I0 =>  inp_feat(115), I1 =>  inp_feat(141), I2 =>  inp_feat(509), I3 =>  inp_feat(273), I4 =>  inp_feat(270), I5 =>  inp_feat(26), I6 =>  inp_feat(485), I7 =>  inp_feat(77)); 
C_33_S_4_L_6_inst : LUT8 generic map(INIT => "0100000000000000000000000000000000000000010000000000000000000000100000001000000000000000000000001000000011001000000000000000000000000000000000000000000010000000101000000000000000000000000000001000000010000000100000000000000010000000110011010000000000000100") port map( O =>C_33_S_4_L_6_out, I0 =>  inp_feat(92), I1 =>  inp_feat(286), I2 =>  inp_feat(9), I3 =>  inp_feat(301), I4 =>  inp_feat(178), I5 =>  inp_feat(53), I6 =>  inp_feat(142), I7 =>  inp_feat(469)); 
C_33_S_4_L_7_inst : LUT8 generic map(INIT => "0100000000000000011100001100000011000000100000001100000011000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000100000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_33_S_4_L_7_out, I0 =>  inp_feat(34), I1 =>  inp_feat(151), I2 =>  inp_feat(160), I3 =>  inp_feat(303), I4 =>  inp_feat(222), I5 =>  inp_feat(382), I6 =>  inp_feat(347), I7 =>  inp_feat(241)); 
C_34_S_0_L_0_inst : LUT8 generic map(INIT => "1111111110100011110010001111101010100010001010101000000010001000111100101011100011110000111111110000000000000000100000001011001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_0_L_0_out, I0 =>  inp_feat(247), I1 =>  inp_feat(286), I2 =>  inp_feat(310), I3 =>  inp_feat(160), I4 =>  inp_feat(180), I5 =>  inp_feat(469), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_34_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111010100111101100000000010101011000000001111101000000000111111111000110011001101000011000000000000000000000000000000000011001010000000000000100000000000000000001000000001000000000000001100100100000000100011100000000000000000000000000000000000000000") port map( O =>C_34_S_0_L_1_out, I0 =>  inp_feat(382), I1 =>  inp_feat(509), I2 =>  inp_feat(494), I3 =>  inp_feat(414), I4 =>  inp_feat(310), I5 =>  inp_feat(430), I6 =>  inp_feat(286), I7 =>  inp_feat(77)); 
C_34_S_0_L_2_inst : LUT8 generic map(INIT => "1111111111101110110000000000000011111011001000000000000000000000111100100000000011000000000000001111100100000000110000000000000011101010111011100100000001000000100000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000") port map( O =>C_34_S_0_L_2_out, I0 =>  inp_feat(145), I1 =>  inp_feat(286), I2 =>  inp_feat(161), I3 =>  inp_feat(273), I4 =>  inp_feat(434), I5 =>  inp_feat(310), I6 =>  inp_feat(303), I7 =>  inp_feat(301)); 
C_34_S_0_L_3_inst : LUT8 generic map(INIT => "1110100011001000111000001000000011001000100000001000000000000000101010001000000010101000000000001010100010000000100010000000000011101111111011111100100000000000110011001000100000000000000000001000000010000000100010000000000010000000100010001000000010001000") port map( O =>C_34_S_0_L_3_out, I0 =>  inp_feat(310), I1 =>  inp_feat(414), I2 =>  inp_feat(142), I3 =>  inp_feat(367), I4 =>  inp_feat(505), I5 =>  inp_feat(509), I6 =>  inp_feat(233), I7 =>  inp_feat(154)); 
C_34_S_0_L_4_inst : LUT8 generic map(INIT => "1111111001110100001010100110000011101100010001001110100011000000101000000010000000001000000000000000000010001000000010000000000000100000000000000010100010100000100000000000000011100000111000000010000000000000001000000010000010000000000000000010000010000000") port map( O =>C_34_S_0_L_4_out, I0 =>  inp_feat(367), I1 =>  inp_feat(344), I2 =>  inp_feat(51), I3 =>  inp_feat(469), I4 =>  inp_feat(26), I5 =>  inp_feat(178), I6 =>  inp_feat(207), I7 =>  inp_feat(450)); 
C_34_S_0_L_5_inst : LUT8 generic map(INIT => "1111110011111010111110001111111111111111100011001000000000000000101000001010000000000000100000001010000000000000101000000000000010111110100010111000100010000000101000100010000000000000000000001000000000000000000000000010000000000000000000000000000000000000") port map( O =>C_34_S_0_L_5_out, I0 =>  inp_feat(48), I1 =>  inp_feat(212), I2 =>  inp_feat(484), I3 =>  inp_feat(301), I4 =>  inp_feat(344), I5 =>  inp_feat(170), I6 =>  inp_feat(382), I7 =>  inp_feat(448)); 
C_34_S_0_L_6_inst : LUT8 generic map(INIT => "1001110011101111110110100000101011011111010111101101000100001100101000001010000011001000100010001100110010001100110110001000110010010000100000001011000000000000000000010100110001011000000000001001000010100000110010001000100000000000000001001101100010001000") port map( O =>C_34_S_0_L_6_out, I0 =>  inp_feat(248), I1 =>  inp_feat(161), I2 =>  inp_feat(171), I3 =>  inp_feat(308), I4 =>  inp_feat(156), I5 =>  inp_feat(180), I6 =>  inp_feat(26), I7 =>  inp_feat(218)); 
C_34_S_0_L_7_inst : LUT8 generic map(INIT => "1110111011001000101010101100010010100010001011111010101010101100110001100000000000000000000000000000000000100111101000001010001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_0_L_7_out, I0 =>  inp_feat(12), I1 =>  inp_feat(344), I2 =>  inp_feat(302), I3 =>  inp_feat(86), I4 =>  inp_feat(427), I5 =>  inp_feat(237), I6 =>  inp_feat(218), I7 =>  inp_feat(257)); 
C_34_S_1_L_0_inst : LUT8 generic map(INIT => "1111111110100011110010001111101010100010001010101000000010001000111100101011100011110000111111110000000000000000100000001011001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_1_L_0_out, I0 =>  inp_feat(247), I1 =>  inp_feat(286), I2 =>  inp_feat(310), I3 =>  inp_feat(160), I4 =>  inp_feat(180), I5 =>  inp_feat(469), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_34_S_1_L_1_inst : LUT8 generic map(INIT => "1111111111010100111101100000000010101011000000001111101000000000111111111000110011001101000011000000000000000000000000000000000011001010000000000000100000000000000000001000000001000000000000001100100100000000100011100000000000000000000000000000000000000000") port map( O =>C_34_S_1_L_1_out, I0 =>  inp_feat(382), I1 =>  inp_feat(509), I2 =>  inp_feat(494), I3 =>  inp_feat(414), I4 =>  inp_feat(310), I5 =>  inp_feat(430), I6 =>  inp_feat(286), I7 =>  inp_feat(77)); 
C_34_S_1_L_2_inst : LUT8 generic map(INIT => "1111110011110101110011010100000010000000000000000000000000000000110011001110110011000000010000001000000000100000000000000000000011001100111000000100000000000000100010001010000000000000000000001110000010100000000000000000000010000000101000000000000000000000") port map( O =>C_34_S_1_L_2_out, I0 =>  inp_feat(351), I1 =>  inp_feat(430), I2 =>  inp_feat(161), I3 =>  inp_feat(41), I4 =>  inp_feat(344), I5 =>  inp_feat(274), I6 =>  inp_feat(485), I7 =>  inp_feat(103)); 
C_34_S_1_L_3_inst : LUT8 generic map(INIT => "1111111111000100111011101000100111111111100010001010111010001000101000001000000010100000000000001010000000000000000000000000000011111011100000001100101100000000111110111100000011111111000000001000000001000000000000000000000011000000110000000000000000000000") port map( O =>C_34_S_1_L_3_out, I0 =>  inp_feat(365), I1 =>  inp_feat(505), I2 =>  inp_feat(425), I3 =>  inp_feat(420), I4 =>  inp_feat(244), I5 =>  inp_feat(154), I6 =>  inp_feat(382), I7 =>  inp_feat(56)); 
C_34_S_1_L_4_inst : LUT8 generic map(INIT => "1110100011001000111100001100000011001010010001000000000000000000101100011010010000110000101000001111110111110101001000000000000011011001010000010011000001110000000100010000000000010000000000000011000100010000001100000001000000010001000100010011000000000001") port map( O =>C_34_S_1_L_4_out, I0 =>  inp_feat(160), I1 =>  inp_feat(204), I2 =>  inp_feat(303), I3 =>  inp_feat(469), I4 =>  inp_feat(301), I5 =>  inp_feat(310), I6 =>  inp_feat(286), I7 =>  inp_feat(142)); 
C_34_S_1_L_5_inst : LUT8 generic map(INIT => "1110110011001000111110101010110011100101100000001111010111000100110011111100000011111001000000001000010100000000111100011000000010101001000010001010101011000000011011011000010011111111111011000000000100000000000000000000000000000000000000000010000000000000") port map( O =>C_34_S_1_L_5_out, I0 =>  inp_feat(347), I1 =>  inp_feat(301), I2 =>  inp_feat(367), I3 =>  inp_feat(303), I4 =>  inp_feat(180), I5 =>  inp_feat(200), I6 =>  inp_feat(386), I7 =>  inp_feat(142)); 
C_34_S_1_L_6_inst : LUT8 generic map(INIT => "1111011111100010111010101010100010001000000000001010101010001000111000100100001000100010100000101000000000000000001000000000000011000000111000001000000000000000100000000000000000000000000000001100000011000000000000000000000000000000000000000010000000000000") port map( O =>C_34_S_1_L_6_out, I0 =>  inp_feat(389), I1 =>  inp_feat(444), I2 =>  inp_feat(367), I3 =>  inp_feat(406), I4 =>  inp_feat(56), I5 =>  inp_feat(303), I6 =>  inp_feat(382), I7 =>  inp_feat(207)); 
C_34_S_1_L_7_inst : LUT8 generic map(INIT => "1110101011111010101010001110100011110000101010111000000000000000101000001010101010000000000000000101110010001000100000000000000011110000111110100100100011001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_1_L_7_out, I0 =>  inp_feat(406), I1 =>  inp_feat(301), I2 =>  inp_feat(310), I3 =>  inp_feat(286), I4 =>  inp_feat(470), I5 =>  inp_feat(344), I6 =>  inp_feat(427), I7 =>  inp_feat(247)); 
C_34_S_2_L_0_inst : LUT8 generic map(INIT => "1111111110100011110010001111101010100010001010101000000010001000111100101011100011110000111111110000000000000000100000001011001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_2_L_0_out, I0 =>  inp_feat(247), I1 =>  inp_feat(286), I2 =>  inp_feat(310), I3 =>  inp_feat(160), I4 =>  inp_feat(180), I5 =>  inp_feat(469), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_34_S_2_L_1_inst : LUT8 generic map(INIT => "1111111111010100111101100000000010101011000000001111101000000000111111111000110011001101000011000000000000000000000000000000000011001010000000000000100000000000000000001000000001000000000000001100100100000000100011100000000000000000000000000000000000000000") port map( O =>C_34_S_2_L_1_out, I0 =>  inp_feat(382), I1 =>  inp_feat(509), I2 =>  inp_feat(494), I3 =>  inp_feat(414), I4 =>  inp_feat(310), I5 =>  inp_feat(430), I6 =>  inp_feat(286), I7 =>  inp_feat(77)); 
C_34_S_2_L_2_inst : LUT8 generic map(INIT => "0000110011001000111111001110010011111010000000000010101000000000111011100100010011101110010000001010101000000000101010100000000011111000111100000100000010000000110010000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_2_L_2_out, I0 =>  inp_feat(156), I1 =>  inp_feat(420), I2 =>  inp_feat(506), I3 =>  inp_feat(326), I4 =>  inp_feat(431), I5 =>  inp_feat(485), I6 =>  inp_feat(215), I7 =>  inp_feat(103)); 
C_34_S_2_L_3_inst : LUT8 generic map(INIT => "1111111110011000100010110000000011100100011100001000000001000000110011001100000011000000010000000000000000000000000000000000000011101100111110000100000011000000100001001100000010000000110100001100110011001000110001001100000000000100100000000000000001000000") port map( O =>C_34_S_2_L_3_out, I0 =>  inp_feat(286), I1 =>  inp_feat(207), I2 =>  inp_feat(170), I3 =>  inp_feat(365), I4 =>  inp_feat(382), I5 =>  inp_feat(310), I6 =>  inp_feat(301), I7 =>  inp_feat(154)); 
C_34_S_2_L_4_inst : LUT8 generic map(INIT => "1110101011001100111010101100100010001010100010000000000000000000110010101000000010000000000000001100101010000010000000000000000011010000100000001111000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_2_L_4_out, I0 =>  inp_feat(158), I1 =>  inp_feat(112), I2 =>  inp_feat(301), I3 =>  inp_feat(319), I4 =>  inp_feat(386), I5 =>  inp_feat(430), I6 =>  inp_feat(77), I7 =>  inp_feat(191)); 
C_34_S_2_L_5_inst : LUT8 generic map(INIT => "1111101011001110111110111000101011101010100010000100001000000000111010101100001011001000000000001000000000000000000000000000000011100000100000001000000000000000000000000000000000000000000000001100000010000000100000000000000000000000000000000000000000000000") port map( O =>C_34_S_2_L_5_out, I0 =>  inp_feat(303), I1 =>  inp_feat(115), I2 =>  inp_feat(301), I3 =>  inp_feat(319), I4 =>  inp_feat(483), I5 =>  inp_feat(386), I6 =>  inp_feat(77), I7 =>  inp_feat(192)); 
C_34_S_2_L_6_inst : LUT8 generic map(INIT => "1100110011000000110100000101000011111100000000000101001000000000110111001101000011010100000100001101110000000000010011000000000011000000100000001100000011110000000000000000000000000000000000001101100011000000110000001000000010000000100000001000000000000000") port map( O =>C_34_S_2_L_6_out, I0 =>  inp_feat(145), I1 =>  inp_feat(430), I2 =>  inp_feat(147), I3 =>  inp_feat(301), I4 =>  inp_feat(448), I5 =>  inp_feat(303), I6 =>  inp_feat(494), I7 =>  inp_feat(92)); 
C_34_S_2_L_7_inst : LUT8 generic map(INIT => "1111111100101101110011001101110001100000100000001100010001001100011000000110000011010000110100000000000000000000000000000000000011111111111101111101000011010000000000000000000001000000000000001111110000011000111100001101000000000000000000000000000000000000") port map( O =>C_34_S_2_L_7_out, I0 =>  inp_feat(178), I1 =>  inp_feat(470), I2 =>  inp_feat(105), I3 =>  inp_feat(303), I4 =>  inp_feat(26), I5 =>  inp_feat(342), I6 =>  inp_feat(509), I7 =>  inp_feat(210)); 
C_34_S_3_L_0_inst : LUT8 generic map(INIT => "1111111110100011110010001111101010100010001010101000000010001000111100101011100011110000111111110000000000000000100000001011001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_3_L_0_out, I0 =>  inp_feat(247), I1 =>  inp_feat(286), I2 =>  inp_feat(310), I3 =>  inp_feat(160), I4 =>  inp_feat(180), I5 =>  inp_feat(469), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_34_S_3_L_1_inst : LUT8 generic map(INIT => "1101111100001000111011110000000011011010000000000000000000000000101010100000000010100000000000000000000000000000000000000000000011101000000000000000000000000000010010000000001000000000000000001010100000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_3_L_1_out, I0 =>  inp_feat(233), I1 =>  inp_feat(301), I2 =>  inp_feat(351), I3 =>  inp_feat(257), I4 =>  inp_feat(264), I5 =>  inp_feat(430), I6 =>  inp_feat(286), I7 =>  inp_feat(77)); 
C_34_S_3_L_2_inst : LUT8 generic map(INIT => "1111101111100010111011100100010011111110110000001010101011001000111110110110001001100000000000000000000001000000000000000000000011101010010010001110101001000000001010101000000000000010000000100100000001000000010000000000000000000000000000000000000000000000") port map( O =>C_34_S_3_L_2_out, I0 =>  inp_feat(156), I1 =>  inp_feat(362), I2 =>  inp_feat(295), I3 =>  inp_feat(218), I4 =>  inp_feat(41), I5 =>  inp_feat(161), I6 =>  inp_feat(48), I7 =>  inp_feat(303)); 
C_34_S_3_L_3_inst : LUT8 generic map(INIT => "1110111010000010111100100000000001101100000010001100000001000100110001000100000001000100000000001100010000000100010001000000000011111110101010001111101011101010110111000000100010001000000010001100110010000000100110000000000011000100000000000000000000000000") port map( O =>C_34_S_3_L_3_out, I0 =>  inp_feat(371), I1 =>  inp_feat(319), I2 =>  inp_feat(373), I3 =>  inp_feat(218), I4 =>  inp_feat(469), I5 =>  inp_feat(310), I6 =>  inp_feat(383), I7 =>  inp_feat(26)); 
C_34_S_3_L_4_inst : LUT8 generic map(INIT => "1011101110100000101000001100000010101000101100001100000010010000110111001100110011010000110100001000100000000000000000000000000010101000101000001010000010100000101000001010000010100000101000001010100000000000000000001000000000100000001000001010000000000000") port map( O =>C_34_S_3_L_4_out, I0 =>  inp_feat(142), I1 =>  inp_feat(212), I2 =>  inp_feat(262), I3 =>  inp_feat(201), I4 =>  inp_feat(172), I5 =>  inp_feat(433), I6 =>  inp_feat(383), I7 =>  inp_feat(495)); 
C_34_S_3_L_5_inst : LUT8 generic map(INIT => "1110111011101000111111101111101011111100001100001010100010100000110000001000000010100010101000001000000000000000100000000000000011111100001100001000000010010000010001001111000000000000100000000100000000000000000000000000000000000000010000000000000000000000") port map( O =>C_34_S_3_L_5_out, I0 =>  inp_feat(31), I1 =>  inp_feat(464), I2 =>  inp_feat(34), I3 =>  inp_feat(301), I4 =>  inp_feat(156), I5 =>  inp_feat(271), I6 =>  inp_feat(77), I7 =>  inp_feat(382)); 
C_34_S_3_L_6_inst : LUT8 generic map(INIT => "1111110011111110111011001110010010000100000011110000110000001100111010001010101011011100000000000000000010001000000001000000000011100000000000001110110010100000000000000000000001000100000000000100000000000000110001000000000000000000000000000100010000000000") port map( O =>C_34_S_3_L_6_out, I0 =>  inp_feat(286), I1 =>  inp_feat(218), I2 =>  inp_feat(367), I3 =>  inp_feat(103), I4 =>  inp_feat(9), I5 =>  inp_feat(227), I6 =>  inp_feat(303), I7 =>  inp_feat(247)); 
C_34_S_3_L_7_inst : LUT8 generic map(INIT => "1101110011111000110111001000000010110000101000000001000000000000100000001100100000000000000010000000000000001000000000000000100011111000100010000100110000000000000000001000100000000000000000000000100010001000000000000000100000000000100010000000000010001000") port map( O =>C_34_S_3_L_7_out, I0 =>  inp_feat(111), I1 =>  inp_feat(310), I2 =>  inp_feat(13), I3 =>  inp_feat(172), I4 =>  inp_feat(247), I5 =>  inp_feat(207), I6 =>  inp_feat(97), I7 =>  inp_feat(358)); 
C_34_S_4_L_0_inst : LUT8 generic map(INIT => "1111111110100011110010001111101010100010001010101000000010001000111100101011100011110000111111110000000000000000100000001011001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_4_L_0_out, I0 =>  inp_feat(247), I1 =>  inp_feat(286), I2 =>  inp_feat(310), I3 =>  inp_feat(160), I4 =>  inp_feat(180), I5 =>  inp_feat(469), I6 =>  inp_feat(142), I7 =>  inp_feat(257)); 
C_34_S_4_L_1_inst : LUT8 generic map(INIT => "1101111100001000111011110000000011011010000000000000000000000000101010100000000010100000000000000000000000000000000000000000000011101000000000000000000000000000010010000000001000000000000000001010100000000000000000000000000000000000000000000000000000000000") port map( O =>C_34_S_4_L_1_out, I0 =>  inp_feat(233), I1 =>  inp_feat(301), I2 =>  inp_feat(351), I3 =>  inp_feat(257), I4 =>  inp_feat(264), I5 =>  inp_feat(430), I6 =>  inp_feat(286), I7 =>  inp_feat(77)); 
C_34_S_4_L_2_inst : LUT8 generic map(INIT => "1111101111100010111011100100010011111110110000001010101011001000111110110110001001100000000000000000000001000000000000000000000011101010010010001110101001000000001010101000000000000010000000100100000001000000010000000000000000000000000000000000000000000000") port map( O =>C_34_S_4_L_2_out, I0 =>  inp_feat(156), I1 =>  inp_feat(362), I2 =>  inp_feat(295), I3 =>  inp_feat(218), I4 =>  inp_feat(41), I5 =>  inp_feat(161), I6 =>  inp_feat(48), I7 =>  inp_feat(303)); 
C_34_S_4_L_3_inst : LUT8 generic map(INIT => "1110111010000010111100100000000001101100000010001100000001000100110001000100000001000100000000001100010000000100010001000000000011111110101010001111101011101010110111000000100010001000000010001100110010000000100110000000000011000100000000000000000000000000") port map( O =>C_34_S_4_L_3_out, I0 =>  inp_feat(371), I1 =>  inp_feat(319), I2 =>  inp_feat(373), I3 =>  inp_feat(218), I4 =>  inp_feat(469), I5 =>  inp_feat(310), I6 =>  inp_feat(383), I7 =>  inp_feat(26)); 
C_34_S_4_L_4_inst : LUT8 generic map(INIT => "1111110011100100110010001100110011100000110111000000000001001100111010001000000000000000100000001000100000000000000000000000000011110000000000001000000000000000000000000000000000000000000000001111000000000000100000000000000000000000000000000000000000000000") port map( O =>C_34_S_4_L_4_out, I0 =>  inp_feat(399), I1 =>  inp_feat(303), I2 =>  inp_feat(239), I3 =>  inp_feat(215), I4 =>  inp_feat(13), I5 =>  inp_feat(147), I6 =>  inp_feat(186), I7 =>  inp_feat(495)); 
C_34_S_4_L_5_inst : LUT8 generic map(INIT => "1111110000111100111100001101000011001100100000001100000001000000111011001110111110101000101000001010000010101000101000001010000001000000000000000000000000000000110000000000000001000000000000001100000010001000001000000000000010000000100000001010000010100000") port map( O =>C_34_S_4_L_5_out, I0 =>  inp_feat(331), I1 =>  inp_feat(186), I2 =>  inp_feat(92), I3 =>  inp_feat(467), I4 =>  inp_feat(319), I5 =>  inp_feat(151), I6 =>  inp_feat(178), I7 =>  inp_feat(77)); 
C_34_S_4_L_6_inst : LUT8 generic map(INIT => "1111111011010100111111001000000011100000111111001000000010100000111111000000000011111100000000001010000010000000000000000010000011001100100001001100110001000000000000000000000000000100000000001000000000000000000010000000000010100000000001000100000000000000") port map( O =>C_34_S_4_L_6_out, I0 =>  inp_feat(382), I1 =>  inp_feat(352), I2 =>  inp_feat(367), I3 =>  inp_feat(406), I4 =>  inp_feat(115), I5 =>  inp_feat(344), I6 =>  inp_feat(310), I7 =>  inp_feat(161)); 
C_34_S_4_L_7_inst : LUT8 generic map(INIT => "1111110111110001110000001111000111001001100000001100000000000000111111011011100000000000011100111000010000000000000000000000000111111101110100000110010011110001000000000000000000000000000100000000110100000000000000000011010000000000100000000000000000000000") port map( O =>C_34_S_4_L_7_out, I0 =>  inp_feat(180), I1 =>  inp_feat(383), I2 =>  inp_feat(303), I3 =>  inp_feat(204), I4 =>  inp_feat(142), I5 =>  inp_feat(207), I6 =>  inp_feat(310), I7 =>  inp_feat(509)); 
C_35_S_0_L_0_inst : LUT8 generic map(INIT => "1111111010101100111011100000101011101110101011001010101010101000110110001010100000000000110000001100110011101100110011000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_0_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(247), I2 =>  inp_feat(229), I3 =>  inp_feat(31), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_35_S_0_L_1_inst : LUT8 generic map(INIT => "1111100111111101101110011001000000001000000000000000000000000000111110011011000100010001000000000000000000000000000000000000000010111000000000000011001100000000000000000000000000000000000000001000100000000000100010000000000000000000000000000000000000000000") port map( O =>C_35_S_0_L_1_out, I0 =>  inp_feat(105), I1 =>  inp_feat(160), I2 =>  inp_feat(218), I3 =>  inp_feat(310), I4 =>  inp_feat(48), I5 =>  inp_feat(257), I6 =>  inp_feat(139), I7 =>  inp_feat(157)); 
C_35_S_0_L_2_inst : LUT8 generic map(INIT => "1010101011000100111011011100100000100010100000001011100100010000000000000000000010000000000000001000000000000001000000000000000011000001110100001011000000010001100100010001000010110011000100011101000111010000000100010001000110010000000100000101000100010101") port map( O =>C_35_S_0_L_2_out, I0 =>  inp_feat(279), I1 =>  inp_feat(314), I2 =>  inp_feat(161), I3 =>  inp_feat(373), I4 =>  inp_feat(286), I5 =>  inp_feat(239), I6 =>  inp_feat(19), I7 =>  inp_feat(154)); 
C_35_S_0_L_3_inst : LUT8 generic map(INIT => "1101100010001000111111101110000011111100100000001111110000000000111010101010000010101010101000000000000000000000001000000000000011101100000000001110110000000000110010000000000011001100000000001110101000000000101010100000000000000000000000001000100000000000") port map( O =>C_35_S_0_L_3_out, I0 =>  inp_feat(218), I1 =>  inp_feat(86), I2 =>  inp_feat(303), I3 =>  inp_feat(193), I4 =>  inp_feat(154), I5 =>  inp_feat(315), I6 =>  inp_feat(120), I7 =>  inp_feat(93)); 
C_35_S_0_L_4_inst : LUT8 generic map(INIT => "1011011111000000110100001100000010110111010000000010000001000000100011001000000000000000100000000100000000000000010000000000000011111010110000000011000000000000111011100100000000100000010000001000000000000000000000000000000011001100000000000000000000000000") port map( O =>C_35_S_0_L_4_out, I0 =>  inp_feat(201), I1 =>  inp_feat(444), I2 =>  inp_feat(48), I3 =>  inp_feat(332), I4 =>  inp_feat(161), I5 =>  inp_feat(469), I6 =>  inp_feat(430), I7 =>  inp_feat(289)); 
C_35_S_0_L_5_inst : LUT8 generic map(INIT => "1111110010111111110011000000000010111000100100001000000000000000111100001010000000010000000000001110000010100000000000000000000000011000000000100000000000000000000100000001100100000000000000000111000010000000001100000000000011110000100000000001000000000000") port map( O =>C_35_S_0_L_5_out, I0 =>  inp_feat(347), I1 =>  inp_feat(90), I2 =>  inp_feat(17), I3 =>  inp_feat(285), I4 =>  inp_feat(470), I5 =>  inp_feat(301), I6 =>  inp_feat(160), I7 =>  inp_feat(142)); 
C_35_S_0_L_6_inst : LUT8 generic map(INIT => "1111101011000000110110000000000011000000110010001100000011000000111000101000000000000000010000001000000010000000110000001000000011011011000000000001001100000000100010001000100011000000100000000000000100001000101000100000000010000000100010000100000010000000") port map( O =>C_35_S_0_L_6_out, I0 =>  inp_feat(448), I1 =>  inp_feat(333), I2 =>  inp_feat(310), I3 =>  inp_feat(227), I4 =>  inp_feat(450), I5 =>  inp_feat(39), I6 =>  inp_feat(469), I7 =>  inp_feat(296)); 
C_35_S_0_L_7_inst : LUT8 generic map(INIT => "1110110011101000111101111000000011101010110010101010000000000000111111111111111111011101111101111010101010101010000000000000000010001000110010001110010000000000100000101100001000000000000000000000001000000010000000000000000000000010000000000000000000000000") port map( O =>C_35_S_0_L_7_out, I0 =>  inp_feat(382), I1 =>  inp_feat(52), I2 =>  inp_feat(509), I3 =>  inp_feat(172), I4 =>  inp_feat(74), I5 =>  inp_feat(432), I6 =>  inp_feat(154), I7 =>  inp_feat(77)); 
C_35_S_1_L_0_inst : LUT8 generic map(INIT => "1111111010101100111011100000101011101110101011001010101010101000110110001010100000000000110000001100110011101100110011000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_1_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(247), I2 =>  inp_feat(229), I3 =>  inp_feat(31), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_35_S_1_L_1_inst : LUT8 generic map(INIT => "1111101011111000111110101111000000000000000000000000000000110000110110001100000011111100101101000000000000000000000000000000000010001000110100001101000000110000000000000000000000000000000000001100100010001100000000000000000000000000000000000000000000000000") port map( O =>C_35_S_1_L_1_out, I0 =>  inp_feat(301), I1 =>  inp_feat(478), I2 =>  inp_feat(303), I3 =>  inp_feat(218), I4 =>  inp_feat(248), I5 =>  inp_feat(257), I6 =>  inp_feat(139), I7 =>  inp_feat(157)); 
C_35_S_1_L_2_inst : LUT8 generic map(INIT => "1111111111010001010011100100110011000000100000001000000010000000111110001111000000000001100001001100000010000000000000000000000011011111100011110000111010001101100000001000000010000000100000001000000011001000000010000000110010000000100000000000000000000000") port map( O =>C_35_S_1_L_2_out, I0 =>  inp_feat(286), I1 =>  inp_feat(310), I2 =>  inp_feat(371), I3 =>  inp_feat(108), I4 =>  inp_feat(509), I5 =>  inp_feat(432), I6 =>  inp_feat(155), I7 =>  inp_feat(154)); 
C_35_S_1_L_3_inst : LUT8 generic map(INIT => "1111111111000000111110111100100011111100110001000000000010000000101000001000000010000000000000000000000010000000000000000000000010110000100000000000000000000000101100001000100000000000000000000000000010001000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_1_L_3_out, I0 =>  inp_feat(19), I1 =>  inp_feat(119), I2 =>  inp_feat(430), I3 =>  inp_feat(478), I4 =>  inp_feat(48), I5 =>  inp_feat(328), I6 =>  inp_feat(466), I7 =>  inp_feat(161)); 
C_35_S_1_L_4_inst : LUT8 generic map(INIT => "1111011011111010111101001110101011001110100000001110000010000000111100101000000011100000000000000111111100000000111100000000000010100000000000001000000010000000101000100000000010000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_1_L_4_out, I0 =>  inp_feat(92), I1 =>  inp_feat(216), I2 =>  inp_feat(310), I3 =>  inp_feat(107), I4 =>  inp_feat(509), I5 =>  inp_feat(201), I6 =>  inp_feat(227), I7 =>  inp_feat(77)); 
C_35_S_1_L_5_inst : LUT8 generic map(INIT => "1111110111101000100000001101000011000000000000000000000000000000110000000001000010000000000000001011000000000000000000000000000011001100111010001110100010110000100000000000000010101000000000000000100000000000010000000000000010000000000000000000000000000000") port map( O =>C_35_S_1_L_5_out, I0 =>  inp_feat(244), I1 =>  inp_feat(112), I2 =>  inp_feat(470), I3 =>  inp_feat(48), I4 =>  inp_feat(5), I5 =>  inp_feat(161), I6 =>  inp_feat(179), I7 =>  inp_feat(171)); 
C_35_S_1_L_6_inst : LUT8 generic map(INIT => "1111111011111100111010001010000011111010000100001000100000000000110010000010000011000000101000001000100000000000000000000000000001011100101011100000000000000000101100000000000000000000000000000000000000101000000000000000000000001000001000000000000000000000") port map( O =>C_35_S_1_L_6_out, I0 =>  inp_feat(303), I1 =>  inp_feat(218), I2 =>  inp_feat(5), I3 =>  inp_feat(448), I4 =>  inp_feat(57), I5 =>  inp_feat(48), I6 =>  inp_feat(112), I7 =>  inp_feat(142)); 
C_35_S_1_L_7_inst : LUT8 generic map(INIT => "1110111011000100111011001100000010100000000000001100000011001000101011000000000000000000000000001010000000000000000000000000000001111100001000000010000010101010000100000000000000000000000000001111111100001000000000000000000000000010000000000000000000000000") port map( O =>C_35_S_1_L_7_out, I0 =>  inp_feat(303), I1 =>  inp_feat(171), I2 =>  inp_feat(509), I3 =>  inp_feat(213), I4 =>  inp_feat(216), I5 =>  inp_feat(207), I6 =>  inp_feat(485), I7 =>  inp_feat(302)); 
C_35_S_2_L_0_inst : LUT8 generic map(INIT => "1111111010101100111011100000101011101110101011001010101010101000110110001010100000000000110000001100110011101100110011000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_2_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(247), I2 =>  inp_feat(229), I3 =>  inp_feat(31), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_35_S_2_L_1_inst : LUT8 generic map(INIT => "1111111011001100111000100000100011111010111011001110101000000001000001000000010000000000000000000000000000000000000000000000000000101100010011001000000000000000111011101100110011000000010000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_2_L_1_out, I0 =>  inp_feat(218), I1 =>  inp_feat(310), I2 =>  inp_feat(248), I3 =>  inp_feat(301), I4 =>  inp_feat(303), I5 =>  inp_feat(154), I6 =>  inp_feat(257), I7 =>  inp_feat(157)); 
C_35_S_2_L_2_inst : LUT8 generic map(INIT => "1111111011110000110010001100000011000000111000001100000011000000000010001000000011001000100000000000000010101000100000001000000010111010111010001000000011000000000000001010000000000000100000001111000111000000000000001000000000000000101000000000000010000000") port map( O =>C_35_S_2_L_2_out, I0 =>  inp_feat(303), I1 =>  inp_feat(218), I2 =>  inp_feat(142), I3 =>  inp_feat(68), I4 =>  inp_feat(205), I5 =>  inp_feat(264), I6 =>  inp_feat(48), I7 =>  inp_feat(432)); 
C_35_S_2_L_3_inst : LUT8 generic map(INIT => "1111111010111011011101100011001110101000101000100000000010111010101000001011000110100000101100110010000000000000001100000010000000000000001100100000000000010000010000000000000000010000000100001100000010110000000000001101000010000000000000000000000000000000") port map( O =>C_35_S_2_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(154), I2 =>  inp_feat(470), I3 =>  inp_feat(56), I4 =>  inp_feat(222), I5 =>  inp_feat(356), I6 =>  inp_feat(351), I7 =>  inp_feat(161)); 
C_35_S_2_L_4_inst : LUT8 generic map(INIT => "1111110011011010100010000000000010100000101010000000000000001000110011001000000000000000000000001000000010001000000000001000000011111100100010001100100010001000100010001000100010000000100010001100110010001000100011001000100010001000100010001000000010001000") port map( O =>C_35_S_2_L_4_out, I0 =>  inp_feat(433), I1 =>  inp_feat(48), I2 =>  inp_feat(53), I3 =>  inp_feat(142), I4 =>  inp_feat(247), I5 =>  inp_feat(451), I6 =>  inp_feat(382), I7 =>  inp_feat(119)); 
C_35_S_2_L_5_inst : LUT8 generic map(INIT => "1111110111001100101111010000000011111000000000001001111100000000111111011000000010011111000000001111000000000000011111110000000011111000000000001111100000000000100010001000000000001000000000001000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_2_L_5_out, I0 =>  inp_feat(347), I1 =>  inp_feat(382), I2 =>  inp_feat(248), I3 =>  inp_feat(48), I4 =>  inp_feat(468), I5 =>  inp_feat(53), I6 =>  inp_feat(485), I7 =>  inp_feat(244)); 
C_35_S_2_L_6_inst : LUT8 generic map(INIT => "1111110111111111100011100000110111101000000001011000111000001101110010000000000010001000000000001000100000000000000000000000000011101100111111001100110001001100000000000001000000001100010001010100110011000000000011000100000000000000000000000000000000000000") port map( O =>C_35_S_2_L_6_out, I0 =>  inp_feat(5), I1 =>  inp_feat(310), I2 =>  inp_feat(56), I3 =>  inp_feat(383), I4 =>  inp_feat(142), I5 =>  inp_feat(161), I6 =>  inp_feat(244), I7 =>  inp_feat(222)); 
C_35_S_2_L_7_inst : LUT8 generic map(INIT => "1100110110110100110101000001110011000100010000000100000010000000110010000000100010010000000001001000000000000000110100000000000011100101111001011101010000000101000001000000000001010100010100001111010100000100111101010111010000100000000000000111000000010000") port map( O =>C_35_S_2_L_7_out, I0 =>  inp_feat(394), I1 =>  inp_feat(469), I2 =>  inp_feat(286), I3 =>  inp_feat(301), I4 =>  inp_feat(509), I5 =>  inp_feat(244), I6 =>  inp_feat(119), I7 =>  inp_feat(154)); 
C_35_S_3_L_0_inst : LUT8 generic map(INIT => "1111111010101100111011100000101011101110101011001010101010101000110110001010100000000000110000001100110011101100110011000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_3_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(247), I2 =>  inp_feat(229), I3 =>  inp_feat(31), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_35_S_3_L_1_inst : LUT8 generic map(INIT => "1111111011001100111000100000100011111010111011001110101000000001000001000000010000000000000000000000000000000000000000000000000000101100010011001000000000000000111011101100110011000000010000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_3_L_1_out, I0 =>  inp_feat(218), I1 =>  inp_feat(310), I2 =>  inp_feat(248), I3 =>  inp_feat(301), I4 =>  inp_feat(303), I5 =>  inp_feat(154), I6 =>  inp_feat(257), I7 =>  inp_feat(157)); 
C_35_S_3_L_2_inst : LUT8 generic map(INIT => "1111111011110000110010001100000011000000111000001100000011000000000010001000000011001000100000000000000010101000100000001000000010111010111010001000000011000000000000001010000000000000100000001111000111000000000000001000000000000000101000000000000010000000") port map( O =>C_35_S_3_L_2_out, I0 =>  inp_feat(303), I1 =>  inp_feat(218), I2 =>  inp_feat(142), I3 =>  inp_feat(68), I4 =>  inp_feat(205), I5 =>  inp_feat(264), I6 =>  inp_feat(48), I7 =>  inp_feat(432)); 
C_35_S_3_L_3_inst : LUT8 generic map(INIT => "1111111011110100110110000101010011110000111100000000000010110100101010101110111010001000110011000000100000000000100010001000010000000000010001000000000000001100000010000000000000001000000001001010101011101110000000000000110000001000000000000000000000000000") port map( O =>C_35_S_3_L_3_out, I0 =>  inp_feat(485), I1 =>  inp_feat(244), I2 =>  inp_feat(331), I3 =>  inp_feat(56), I4 =>  inp_feat(222), I5 =>  inp_feat(356), I6 =>  inp_feat(351), I7 =>  inp_feat(161)); 
C_35_S_3_L_4_inst : LUT8 generic map(INIT => "1111100011111010111011000000000011111001000000001110100000000000110000001100100011001000010000001100100000000000110010000000000011111010101110100000000000000000000000000000000000001000000000001100101011001000100010000100100010001000000010001000110000001000") port map( O =>C_35_S_3_L_4_out, I0 =>  inp_feat(376), I1 =>  inp_feat(391), I2 =>  inp_feat(142), I3 =>  inp_feat(31), I4 =>  inp_feat(5), I5 =>  inp_feat(354), I6 =>  inp_feat(286), I7 =>  inp_feat(53)); 
C_35_S_3_L_5_inst : LUT8 generic map(INIT => "1111101001001010101010000000000011111000100110001111000000000000111110110100101010000000000000001101100010001000000000000000000011100010100000001110100000000000110000001000000010100000000000000000001100000000000100000000000000000000000000000000000000000000") port map( O =>C_35_S_3_L_5_out, I0 =>  inp_feat(77), I1 =>  inp_feat(448), I2 =>  inp_feat(92), I3 =>  inp_feat(382), I4 =>  inp_feat(242), I5 =>  inp_feat(303), I6 =>  inp_feat(53), I7 =>  inp_feat(244)); 
C_35_S_3_L_6_inst : LUT8 generic map(INIT => "1111101010101000110101100000000011011001000000000101010110000000101011000000000000000000000000001000100000000000000000000000000011111111101110011111111110100000101110011010100010111111101101100010111100000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_3_L_6_out, I0 =>  inp_feat(301), I1 =>  inp_feat(367), I2 =>  inp_feat(509), I3 =>  inp_feat(310), I4 =>  inp_feat(451), I5 =>  inp_feat(382), I6 =>  inp_feat(244), I7 =>  inp_feat(154)); 
C_35_S_3_L_7_inst : LUT8 generic map(INIT => "1111110110111011101010100000001011110000000000001000000000000000111111101010100010101000000000001101110010000100100010000000000011101011101100111000100010000000111000001100000010000000000000001110000000100000100000000000000010000000000000001000000000000000") port map( O =>C_35_S_3_L_7_out, I0 =>  inp_feat(48), I1 =>  inp_feat(357), I2 =>  inp_feat(372), I3 =>  inp_feat(301), I4 =>  inp_feat(468), I5 =>  inp_feat(244), I6 =>  inp_feat(201), I7 =>  inp_feat(107)); 
C_35_S_4_L_0_inst : LUT8 generic map(INIT => "1111111010101100111011100000101011101110101011001010101010101000110110001010100000000000110000001100110011101100110011000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_4_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(247), I2 =>  inp_feat(229), I3 =>  inp_feat(31), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_35_S_4_L_1_inst : LUT8 generic map(INIT => "1111111011001100111000100000100011111010111011001110101000000001000001000000010000000000000000000000000000000000000000000000000000101100010011001000000000000000111011101100110011000000010000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_35_S_4_L_1_out, I0 =>  inp_feat(218), I1 =>  inp_feat(310), I2 =>  inp_feat(248), I3 =>  inp_feat(301), I4 =>  inp_feat(303), I5 =>  inp_feat(154), I6 =>  inp_feat(257), I7 =>  inp_feat(157)); 
C_35_S_4_L_2_inst : LUT8 generic map(INIT => "1111111011110000110010001100000011000000111000001100000011000000000010001000000011001000100000000000000010101000100000001000000010111010111010001000000011000000000000001010000000000000100000001111000111000000000000001000000000000000101000000000000010000000") port map( O =>C_35_S_4_L_2_out, I0 =>  inp_feat(303), I1 =>  inp_feat(218), I2 =>  inp_feat(142), I3 =>  inp_feat(68), I4 =>  inp_feat(205), I5 =>  inp_feat(264), I6 =>  inp_feat(48), I7 =>  inp_feat(432)); 
C_35_S_4_L_3_inst : LUT8 generic map(INIT => "1111111011110100110110000101010011110000111100000000000010110100101010101110111010001000110011000000100000000000100010001000010000000000010001000000000000001100000010000000000000001000000001001010101011101110000000000000110000001000000000000000000000000000") port map( O =>C_35_S_4_L_3_out, I0 =>  inp_feat(485), I1 =>  inp_feat(244), I2 =>  inp_feat(331), I3 =>  inp_feat(56), I4 =>  inp_feat(222), I5 =>  inp_feat(356), I6 =>  inp_feat(351), I7 =>  inp_feat(161)); 
C_35_S_4_L_4_inst : LUT8 generic map(INIT => "1111100011110110101110000000000010111011000000001010110000000000110000001100010010000100100000001100010000000000110011000000000011100110111001000000000000000000000000000000000000000100000000001000010111000100010001001000010001001100000001001100110000000100") port map( O =>C_35_S_4_L_4_out, I0 =>  inp_feat(210), I1 =>  inp_feat(391), I2 =>  inp_feat(142), I3 =>  inp_feat(31), I4 =>  inp_feat(5), I5 =>  inp_feat(354), I6 =>  inp_feat(286), I7 =>  inp_feat(53)); 
C_35_S_4_L_5_inst : LUT8 generic map(INIT => "1111101001001010101010000000000011111000100110001111000000000000111110110100101010000000000000001101100010001000000000000000000011100010100000001110100000000000110000001000000010100000000000000000001100000000000100000000000000000000000000000000000000000000") port map( O =>C_35_S_4_L_5_out, I0 =>  inp_feat(77), I1 =>  inp_feat(448), I2 =>  inp_feat(92), I3 =>  inp_feat(382), I4 =>  inp_feat(242), I5 =>  inp_feat(303), I6 =>  inp_feat(53), I7 =>  inp_feat(244)); 
C_35_S_4_L_6_inst : LUT8 generic map(INIT => "1111101011110000101010001100000010110000010000001010100010100000100000000100000010100000000000001010000000000000101000000000000011111111110000001110100011101100101000101110000011100000111100001110100000000000000010000000000000000000000000000000000000000000") port map( O =>C_35_S_4_L_6_out, I0 =>  inp_feat(448), I1 =>  inp_feat(303), I2 =>  inp_feat(86), I3 =>  inp_feat(53), I4 =>  inp_feat(347), I5 =>  inp_feat(382), I6 =>  inp_feat(244), I7 =>  inp_feat(154)); 
C_35_S_4_L_7_inst : LUT8 generic map(INIT => "1110111111011000111110101101000011001001110000001000000001010000110111101000101010001010000000001000100010000000000000000000000011111010110000001111101011010000000000000000000001100000010100000001101000000000101110100000000000000000000000000000000000010000") port map( O =>C_35_S_4_L_7_out, I0 =>  inp_feat(53), I1 =>  inp_feat(52), I2 =>  inp_feat(154), I3 =>  inp_feat(215), I4 =>  inp_feat(399), I5 =>  inp_feat(321), I6 =>  inp_feat(212), I7 =>  inp_feat(412)); 
C_36_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000001000000000001011101010000010100000000000000000000000001000000000000000000000001010000000000000000000000000000000000000000000000010000000000000101010100000000000000000000000000000000000000000") port map( O =>C_36_S_0_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(141), I2 =>  inp_feat(470), I3 =>  inp_feat(58), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_36_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000100000101000000000000000100000000000000010000000000000000000110010000000000000000010100000001000100010001000000000000000000010001000001010") port map( O =>C_36_S_0_L_1_out, I0 =>  inp_feat(286), I1 =>  inp_feat(218), I2 =>  inp_feat(391), I3 =>  inp_feat(274), I4 =>  inp_feat(382), I5 =>  inp_feat(247), I6 =>  inp_feat(386), I7 =>  inp_feat(77)); 
C_36_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000100010000001100000010000000110000000000000000000000100000001000000000000000000000000000000010000000") port map( O =>C_36_S_0_L_2_out, I0 =>  inp_feat(74), I1 =>  inp_feat(286), I2 =>  inp_feat(178), I3 =>  inp_feat(420), I4 =>  inp_feat(218), I5 =>  inp_feat(161), I6 =>  inp_feat(464), I7 =>  inp_feat(509)); 
C_36_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000010000000000011001000000000000000000000000000100010000000010000001000000000101000100000000000000000000000000010001000000000000000000000001010000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000") port map( O =>C_36_S_0_L_3_out, I0 =>  inp_feat(145), I1 =>  inp_feat(382), I2 =>  inp_feat(472), I3 =>  inp_feat(48), I4 =>  inp_feat(509), I5 =>  inp_feat(403), I6 =>  inp_feat(428), I7 =>  inp_feat(220)); 
C_36_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000000000000000101000000000000010000000110010001000000000000000000000000000000000000000000000000000000010000000101000000010000000100010001111101010000000000000001000001000101010000000000000000") port map( O =>C_36_S_0_L_4_out, I0 =>  inp_feat(382), I1 =>  inp_feat(358), I2 =>  inp_feat(86), I3 =>  inp_feat(77), I4 =>  inp_feat(82), I5 =>  inp_feat(212), I6 =>  inp_feat(448), I7 =>  inp_feat(469)); 
C_36_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000011001000000000000000000000000000000000000000000000101000000000000010110000000000000000000000000000000000000001000000000000000001100011000000000000100000000000000010000000100000001110000000000000111100001000") port map( O =>C_36_S_0_L_5_out, I0 =>  inp_feat(13), I1 =>  inp_feat(136), I2 =>  inp_feat(382), I3 =>  inp_feat(351), I4 =>  inp_feat(222), I5 =>  inp_feat(77), I6 =>  inp_feat(303), I7 =>  inp_feat(301)); 
C_36_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000011001000000000000000000000000000000000000000000000101000000000000010110000000000000000000000000000000000000001000000000000000001100011000000000000100000000000000010000000100000001110000000000000111100001000") port map( O =>C_36_S_0_L_6_out, I0 =>  inp_feat(13), I1 =>  inp_feat(136), I2 =>  inp_feat(382), I3 =>  inp_feat(351), I4 =>  inp_feat(222), I5 =>  inp_feat(77), I6 =>  inp_feat(303), I7 =>  inp_feat(301)); 
C_36_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000011001000000000000000000000000000000000000000000000101000000000000010110000000000000000000000000000000000000001000000000000000001100011000000000000100000000000000010000000100000001110000000000000111100001000") port map( O =>C_36_S_0_L_7_out, I0 =>  inp_feat(13), I1 =>  inp_feat(136), I2 =>  inp_feat(382), I3 =>  inp_feat(351), I4 =>  inp_feat(222), I5 =>  inp_feat(77), I6 =>  inp_feat(303), I7 =>  inp_feat(301)); 
C_36_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000001000000000001011101010000010100000000000000000000000001000000000000000000000001010000000000000000000000000000000000000000000000010000000000000101010100000000000000000000000000000000000000000") port map( O =>C_36_S_1_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(141), I2 =>  inp_feat(470), I3 =>  inp_feat(58), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_36_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000100000000000000000000000000000000000000000000000000000001000100000000000000010000000000010001000100000000000100010001000100010000000000000000000") port map( O =>C_36_S_1_L_1_out, I0 =>  inp_feat(178), I1 =>  inp_feat(58), I2 =>  inp_feat(5), I3 =>  inp_feat(448), I4 =>  inp_feat(331), I5 =>  inp_feat(382), I6 =>  inp_feat(509), I7 =>  inp_feat(77)); 
C_36_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000001000000000000000000000000000100010001000101101000000000000001100100000000000000000011000000111000001110000") port map( O =>C_36_S_1_L_2_out, I0 =>  inp_feat(141), I1 =>  inp_feat(222), I2 =>  inp_feat(262), I3 =>  inp_feat(297), I4 =>  inp_feat(77), I5 =>  inp_feat(358), I6 =>  inp_feat(310), I7 =>  inp_feat(509)); 
C_36_S_1_L_3_inst : LUT8 generic map(INIT => "0000000100011011001100011001111100000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_1_L_3_out, I0 =>  inp_feat(435), I1 =>  inp_feat(142), I2 =>  inp_feat(386), I3 =>  inp_feat(77), I4 =>  inp_feat(407), I5 =>  inp_feat(58), I6 =>  inp_feat(20), I7 =>  inp_feat(390)); 
C_36_S_1_L_4_inst : LUT8 generic map(INIT => "0000000001010001000100000111000000000000000100000101000011010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_1_L_4_out, I0 =>  inp_feat(509), I1 =>  inp_feat(239), I2 =>  inp_feat(178), I3 =>  inp_feat(303), I4 =>  inp_feat(211), I5 =>  inp_feat(430), I6 =>  inp_feat(286), I7 =>  inp_feat(240)); 
C_36_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000100000000010000000100000011000101010100000100010000000101010000010100000000000000000000000000000000000000000000000000000100000000000") port map( O =>C_36_S_1_L_5_out, I0 =>  inp_feat(178), I1 =>  inp_feat(298), I2 =>  inp_feat(303), I3 =>  inp_feat(247), I4 =>  inp_feat(310), I5 =>  inp_feat(367), I6 =>  inp_feat(160), I7 =>  inp_feat(218)); 
C_36_S_1_L_6_inst : LUT8 generic map(INIT => "0000010100001000000000010000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000010011001000000001011111110000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000") port map( O =>C_36_S_1_L_6_out, I0 =>  inp_feat(72), I1 =>  inp_feat(77), I2 =>  inp_feat(247), I3 =>  inp_feat(374), I4 =>  inp_feat(469), I5 =>  inp_feat(248), I6 =>  inp_feat(216), I7 =>  inp_feat(218)); 
C_36_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000010000100010000000000000010000000100000010000000000000000100101000100000000000000000000000000001011000000000000000000000000000000000000000000000000000101010001011100000100000000000000010100000001") port map( O =>C_36_S_1_L_7_out, I0 =>  inp_feat(222), I1 =>  inp_feat(310), I2 =>  inp_feat(448), I3 =>  inp_feat(247), I4 =>  inp_feat(382), I5 =>  inp_feat(344), I6 =>  inp_feat(509), I7 =>  inp_feat(358)); 
C_36_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000001000000000001011101010000010100000000000000000000000001000000000000000000000001010000000000000000000000000000000000000000000000010000000000000101010100000000000000000000000000000000000000000") port map( O =>C_36_S_2_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(141), I2 =>  inp_feat(470), I3 =>  inp_feat(58), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_36_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000100000000000000000000000000000000000000000000000000000001000100000000000000010000000000010001000100000000000100010001000100010000000000000000000") port map( O =>C_36_S_2_L_1_out, I0 =>  inp_feat(178), I1 =>  inp_feat(58), I2 =>  inp_feat(5), I3 =>  inp_feat(448), I4 =>  inp_feat(331), I5 =>  inp_feat(382), I6 =>  inp_feat(509), I7 =>  inp_feat(77)); 
C_36_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000001000000000000000000000000000100010001000101101000000000000001100100000000000000000011000000111000001110000") port map( O =>C_36_S_2_L_2_out, I0 =>  inp_feat(141), I1 =>  inp_feat(222), I2 =>  inp_feat(262), I3 =>  inp_feat(297), I4 =>  inp_feat(77), I5 =>  inp_feat(358), I6 =>  inp_feat(310), I7 =>  inp_feat(509)); 
C_36_S_2_L_3_inst : LUT8 generic map(INIT => "0000000100000000000110010001000000000001000000000000000100000000000000000000000000010011000100000000000100000000001100110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000") port map( O =>C_36_S_2_L_3_out, I0 =>  inp_feat(448), I1 =>  inp_feat(382), I2 =>  inp_feat(77), I3 =>  inp_feat(160), I4 =>  inp_feat(407), I5 =>  inp_feat(186), I6 =>  inp_feat(182), I7 =>  inp_feat(390)); 
C_36_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000100100000000000000000000000000000001000000000001000100000000000000010000000000000000000000000000000000000000000000000000000010011001010000000000000000000000000000010000100110000001100100011001000110000000000000000000000000000000000") port map( O =>C_36_S_2_L_4_out, I0 =>  inp_feat(5), I1 =>  inp_feat(178), I2 =>  inp_feat(448), I3 =>  inp_feat(239), I4 =>  inp_feat(303), I5 =>  inp_feat(261), I6 =>  inp_feat(157), I7 =>  inp_feat(469)); 
C_36_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000001010000000000000000000000000001010101010101000000000100000000000110000000000000000000000000000001000000000100000000000001010") port map( O =>C_36_S_2_L_5_out, I0 =>  inp_feat(178), I1 =>  inp_feat(189), I2 =>  inp_feat(509), I3 =>  inp_feat(105), I4 =>  inp_feat(275), I5 =>  inp_feat(161), I6 =>  inp_feat(177), I7 =>  inp_feat(218)); 
C_36_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000101001001010000000000000000001100100001010100000000000000000000001100000101010001010000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000010000000000000000000000100") port map( O =>C_36_S_2_L_6_out, I0 =>  inp_feat(382), I1 =>  inp_feat(77), I2 =>  inp_feat(161), I3 =>  inp_feat(323), I4 =>  inp_feat(238), I5 =>  inp_feat(239), I6 =>  inp_feat(469), I7 =>  inp_feat(331)); 
C_36_S_2_L_7_inst : LUT8 generic map(INIT => "0001000000010000000000000010000001110000011000000001000001000000001100001010000000110000000100000011000000000000011100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_2_L_7_out, I0 =>  inp_feat(229), I1 =>  inp_feat(161), I2 =>  inp_feat(135), I3 =>  inp_feat(74), I4 =>  inp_feat(373), I5 =>  inp_feat(201), I6 =>  inp_feat(414), I7 =>  inp_feat(286)); 
C_36_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000001000000000001011101010000010100000000000000000000000001000000000000000000000001010000000000000000000000000000000000000000000000010000000000000101010100000000000000000000000000000000000000000") port map( O =>C_36_S_3_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(141), I2 =>  inp_feat(470), I3 =>  inp_feat(58), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_36_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000100000000000000000000000000000000000000000000000000000001000100000000000000010000000000010001000100000000000100010001000100010000000000000000000") port map( O =>C_36_S_3_L_1_out, I0 =>  inp_feat(178), I1 =>  inp_feat(58), I2 =>  inp_feat(5), I3 =>  inp_feat(448), I4 =>  inp_feat(331), I5 =>  inp_feat(382), I6 =>  inp_feat(509), I7 =>  inp_feat(77)); 
C_36_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000001000000000000000000000000000100010001000101101000000000000001100100000000000000000011000000111000001110000") port map( O =>C_36_S_3_L_2_out, I0 =>  inp_feat(141), I1 =>  inp_feat(222), I2 =>  inp_feat(262), I3 =>  inp_feat(297), I4 =>  inp_feat(77), I5 =>  inp_feat(358), I6 =>  inp_feat(310), I7 =>  inp_feat(509)); 
C_36_S_3_L_3_inst : LUT8 generic map(INIT => "0001000001010000111100000011000000110001001100000000000000010000000000000000000000000000000100000000000000010000001100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_3_L_3_out, I0 =>  inp_feat(224), I1 =>  inp_feat(142), I2 =>  inp_feat(351), I3 =>  inp_feat(257), I4 =>  inp_feat(407), I5 =>  inp_feat(186), I6 =>  inp_feat(182), I7 =>  inp_feat(390)); 
C_36_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000100000000100000100001101000000010010010100000000010001110000000000000000000001010000110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_3_L_4_out, I0 =>  inp_feat(448), I1 =>  inp_feat(344), I2 =>  inp_feat(420), I3 =>  inp_feat(161), I4 =>  inp_feat(77), I5 =>  inp_feat(157), I6 =>  inp_feat(303), I7 =>  inp_feat(120)); 
C_36_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000001010000000000000000000000000000000000000000000000010001000000000001000100000000000000010000000100000000000000010000000000000000001101010000000000000000000000000000000110000001000100010000000000011001000000000") port map( O =>C_36_S_3_L_5_out, I0 =>  inp_feat(464), I1 =>  inp_feat(382), I2 =>  inp_feat(475), I3 =>  inp_feat(368), I4 =>  inp_feat(494), I5 =>  inp_feat(48), I6 =>  inp_feat(414), I7 =>  inp_feat(301)); 
C_36_S_3_L_6_inst : LUT8 generic map(INIT => "0000001000001011000000100011001100000000000000000000001000101010010100000000101011110001001110100000000100000000000000000010100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_3_L_6_out, I0 =>  inp_feat(470), I1 =>  inp_feat(247), I2 =>  inp_feat(227), I3 =>  inp_feat(77), I4 =>  inp_feat(469), I5 =>  inp_feat(5), I6 =>  inp_feat(226), I7 =>  inp_feat(286)); 
C_36_S_3_L_7_inst : LUT8 generic map(INIT => "0000000001000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000011100000101000000000010010100001111000000000000000100000000000000000000010000000000000001000000000000000000000000000000") port map( O =>C_36_S_3_L_7_out, I0 =>  inp_feat(61), I1 =>  inp_feat(88), I2 =>  inp_feat(286), I3 =>  inp_feat(303), I4 =>  inp_feat(147), I5 =>  inp_feat(301), I6 =>  inp_feat(235), I7 =>  inp_feat(218)); 
C_36_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000001000000000001011101010000010100000000000000000000000001000000000000000000000001010000000000000000000000000000000000000000000000010000000000000101010100000000000000000000000000000000000000000") port map( O =>C_36_S_4_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(141), I2 =>  inp_feat(470), I3 =>  inp_feat(58), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_36_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000100000000000000000000000000000000000000000000000000000001000100000000000000010000000000010001000100000000000100010001000100010000000000000000000") port map( O =>C_36_S_4_L_1_out, I0 =>  inp_feat(178), I1 =>  inp_feat(58), I2 =>  inp_feat(5), I3 =>  inp_feat(448), I4 =>  inp_feat(331), I5 =>  inp_feat(382), I6 =>  inp_feat(509), I7 =>  inp_feat(77)); 
C_36_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000001000000000000000000000000000100010001000101101000000000000001100100000000000000000011000000111000001110000") port map( O =>C_36_S_4_L_2_out, I0 =>  inp_feat(141), I1 =>  inp_feat(222), I2 =>  inp_feat(262), I3 =>  inp_feat(297), I4 =>  inp_feat(77), I5 =>  inp_feat(358), I6 =>  inp_feat(310), I7 =>  inp_feat(509)); 
C_36_S_4_L_3_inst : LUT8 generic map(INIT => "0001000001010000111100000011000000110001001100000000000000010000000000000000000000000000000100000000000000010000001100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_4_L_3_out, I0 =>  inp_feat(224), I1 =>  inp_feat(142), I2 =>  inp_feat(351), I3 =>  inp_feat(257), I4 =>  inp_feat(407), I5 =>  inp_feat(186), I6 =>  inp_feat(182), I7 =>  inp_feat(390)); 
C_36_S_4_L_4_inst : LUT8 generic map(INIT => "0001000100001010000000000000000000100001001100000000000000000000010000000001100100000000000000000000000101110001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_36_S_4_L_4_out, I0 =>  inp_feat(298), I1 =>  inp_feat(77), I2 =>  inp_feat(475), I3 =>  inp_feat(303), I4 =>  inp_feat(385), I5 =>  inp_feat(450), I6 =>  inp_feat(414), I7 =>  inp_feat(120)); 
C_36_S_4_L_5_inst : LUT8 generic map(INIT => "0000001000000000000000000000000000000010000000000000000000000000000010110000010000000000000000000010101000000000000000000000000000001010000000000000000000000000001010100000000000000001000000000010101000000000000000000000000000101010001000100000000000000000") port map( O =>C_36_S_4_L_5_out, I0 =>  inp_feat(180), I1 =>  inp_feat(435), I2 =>  inp_feat(469), I3 =>  inp_feat(347), I4 =>  inp_feat(237), I5 =>  inp_feat(372), I6 =>  inp_feat(53), I7 =>  inp_feat(414)); 
C_36_S_4_L_6_inst : LUT8 generic map(INIT => "0001000000000000000100000011000000010000000100000000000000000000000000000000000000010000001100000000000000000000000000000101000011010000010100000001000011111000000000000000000001000000000001000000000000000000000100000011000000000000000000000000000000010001") port map( O =>C_36_S_4_L_6_out, I0 =>  inp_feat(218), I1 =>  inp_feat(43), I2 =>  inp_feat(180), I3 =>  inp_feat(373), I4 =>  inp_feat(247), I5 =>  inp_feat(5), I6 =>  inp_feat(291), I7 =>  inp_feat(301)); 
C_36_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000100000001000000010000000000000010000000010000000000000010000001000000011100000000000000100000110100000010001000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000001000000000000") port map( O =>C_36_S_4_L_7_out, I0 =>  inp_feat(373), I1 =>  inp_feat(222), I2 =>  inp_feat(216), I3 =>  inp_feat(77), I4 =>  inp_feat(310), I5 =>  inp_feat(367), I6 =>  inp_feat(448), I7 =>  inp_feat(20)); 
C_37_S_0_L_0_inst : LUT8 generic map(INIT => "1111001111110101111000100000100011110011101010101000000010101010111101111111011100000000010000001111011110101010000000001010101000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_0_L_0_out, I0 =>  inp_feat(286), I1 =>  inp_feat(154), I2 =>  inp_feat(52), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_37_S_0_L_1_inst : LUT8 generic map(INIT => "1111101011101110111000101010001011110010100000000000000000000000110010101100000011000010110000101000001010000000000000000000000000110010110011000000001000000000111100111100100000000000000000001011101011000000000000000100000010110011100000000000000000000000") port map( O =>C_37_S_0_L_1_out, I0 =>  inp_feat(303), I1 =>  inp_feat(314), I2 =>  inp_feat(161), I3 =>  inp_feat(216), I4 =>  inp_feat(435), I5 =>  inp_feat(289), I6 =>  inp_feat(115), I7 =>  inp_feat(365)); 
C_37_S_0_L_2_inst : LUT8 generic map(INIT => "1101111110100000101010101000100111110011111100010000000000001000111010101010100011111000100010001010000010100000000000000000000011001000101000001100000000000000111000000000000000000000000000001101110000000000110100001000000000000000000000000000000000000000") port map( O =>C_37_S_0_L_2_out, I0 =>  inp_feat(303), I1 =>  inp_feat(509), I2 =>  inp_feat(218), I3 =>  inp_feat(406), I4 =>  inp_feat(10), I5 =>  inp_feat(485), I6 =>  inp_feat(31), I7 =>  inp_feat(310)); 
C_37_S_0_L_3_inst : LUT8 generic map(INIT => "1111011111110111111011000000000101111111101111110000110100110110101000001010000010100000100000001000000010000000000000000000000011100000000001000010000000000000001000100000010000000000000000001000000010000000101000001000000000000000000000001000000010000000") port map( O =>C_37_S_0_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(119), I2 =>  inp_feat(347), I3 =>  inp_feat(74), I4 =>  inp_feat(469), I5 =>  inp_feat(382), I6 =>  inp_feat(26), I7 =>  inp_feat(77)); 
C_37_S_0_L_4_inst : LUT8 generic map(INIT => "1110111011101100110011001100110011101110111000001110110001100000111011101110010011101111111010000010000000000000000000000000000010001110111000000000100000000000110000000000000000000000000000001000100010100000001011101010000000000000000000000000000000100000") port map( O =>C_37_S_0_L_4_out, I0 =>  inp_feat(301), I1 =>  inp_feat(303), I2 =>  inp_feat(212), I3 =>  inp_feat(480), I4 =>  inp_feat(469), I5 =>  inp_feat(382), I6 =>  inp_feat(26), I7 =>  inp_feat(77)); 
C_37_S_0_L_5_inst : LUT8 generic map(INIT => "1111111111101110101000001010101011000100110011000000000010000000110010001000000000000000000000001000000010000000100000000000000011111011101000000000000000100010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_0_L_5_out, I0 =>  inp_feat(347), I1 =>  inp_feat(151), I2 =>  inp_feat(142), I3 =>  inp_feat(178), I4 =>  inp_feat(430), I5 =>  inp_feat(161), I6 =>  inp_feat(466), I7 =>  inp_feat(48)); 
C_37_S_0_L_6_inst : LUT8 generic map(INIT => "1111110010001000111011101010001010100000000000001010111010101000111011001000110011101111001000000100000000000000111011110000000011100100111010001010000010001000101000001010000000100000101010101010000011101110101010001000100000000000000000000000000000000000") port map( O =>C_37_S_0_L_6_out, I0 =>  inp_feat(367), I1 =>  inp_feat(218), I2 =>  inp_feat(469), I3 =>  inp_feat(23), I4 =>  inp_feat(26), I5 =>  inp_feat(450), I6 =>  inp_feat(212), I7 =>  inp_feat(331)); 
C_37_S_0_L_7_inst : LUT8 generic map(INIT => "1111110011101000111110001000100011101010001000001000000000000000110000001000000010000000000000001010101000100010111011000000001011111000111110000000000000000000100000001000100010000000100010001010000010110000000000000000000000000000000100000000000000000000") port map( O =>C_37_S_0_L_7_out, I0 =>  inp_feat(382), I1 =>  inp_feat(247), I2 =>  inp_feat(37), I3 =>  inp_feat(52), I4 =>  inp_feat(77), I5 =>  inp_feat(452), I6 =>  inp_feat(480), I7 =>  inp_feat(115)); 
C_37_S_1_L_0_inst : LUT8 generic map(INIT => "1111001111110101111000100000100011110011101010101000000010101010111101111111011100000000010000001111011110101010000000001010101000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_1_L_0_out, I0 =>  inp_feat(286), I1 =>  inp_feat(154), I2 =>  inp_feat(52), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_37_S_1_L_1_inst : LUT8 generic map(INIT => "1111000011100000111100001110100011100000110000001010000010000000111100001100000000000000101100001010000011000000101000000000000000000000101000000000000010000010000000001000000010000000100000000000000010010000000000001000000000000000000000001000000010000000") port map( O =>C_37_S_1_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(301), I2 =>  inp_feat(257), I3 =>  inp_feat(178), I4 =>  inp_feat(364), I5 =>  inp_feat(62), I6 =>  inp_feat(373), I7 =>  inp_feat(430)); 
C_37_S_1_L_2_inst : LUT8 generic map(INIT => "1111000011100010001000001100101010001100110010100000000010101010101000001010001010000000110000101000000010100010100000001000001011101000100000000000000011000000100010001000000000000000000000001000000000000000000000001100000000000000000000000000000000000000") port map( O =>C_37_S_1_L_2_out, I0 =>  inp_feat(77), I1 =>  inp_feat(347), I2 =>  inp_feat(39), I3 =>  inp_feat(216), I4 =>  inp_feat(310), I5 =>  inp_feat(211), I6 =>  inp_feat(424), I7 =>  inp_feat(280)); 
C_37_S_1_L_3_inst : LUT8 generic map(INIT => "1110111011101000111010101110000010100000101000000000000010100000111010000110000010001110101000001001000010100000000000001010000011001100111000001100000011000000000000000010000000000100000000001000010000000000000000001000000000000000000000000000000000000000") port map( O =>C_37_S_1_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(107), I2 =>  inp_feat(466), I3 =>  inp_feat(328), I4 =>  inp_feat(382), I5 =>  inp_feat(430), I6 =>  inp_feat(509), I7 =>  inp_feat(161)); 
C_37_S_1_L_4_inst : LUT8 generic map(INIT => "1111111111111011110101000100010011101011100010111101010000000000000000001000000010001100000000000000000000000000000011000000000010111111110011001111110101000100000000000000000011110000000000001010101010000000111111010000000000000000000000001101110000000000") port map( O =>C_37_S_1_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(303), I2 =>  inp_feat(238), I3 =>  inp_feat(357), I4 =>  inp_feat(9), I5 =>  inp_feat(161), I6 =>  inp_feat(475), I7 =>  inp_feat(390)); 
C_37_S_1_L_5_inst : LUT8 generic map(INIT => "1111101011011010111110000000100011101000000010001010100000000000111010001100100001001000110000000000100000000000000000000000000011001010110010100000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_1_L_5_out, I0 =>  inp_feat(276), I1 =>  inp_feat(13), I2 =>  inp_feat(160), I3 =>  inp_feat(323), I4 =>  inp_feat(364), I5 =>  inp_feat(161), I6 =>  inp_feat(470), I7 =>  inp_feat(48)); 
C_37_S_1_L_6_inst : LUT8 generic map(INIT => "1110100011101000110001000000000011110010010100100100000000000000110011001000100001000100000000001000100000000000000000000000000010101010001010101110000000101000101000100010001000000000001000101000100010000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_1_L_6_out, I0 =>  inp_feat(314), I1 =>  inp_feat(237), I2 =>  inp_feat(373), I3 =>  inp_feat(48), I4 =>  inp_feat(142), I5 =>  inp_feat(376), I6 =>  inp_feat(166), I7 =>  inp_feat(406)); 
C_37_S_1_L_7_inst : LUT8 generic map(INIT => "1110111100001000111100001000001011111111000000001101000000000000111011111000110011110100010001000000111100000000000000000000000011000000000000000010100000001000100010000000000010000000000010001100110010001100111100001111111000000000000000000000000000000000") port map( O =>C_37_S_1_L_7_out, I0 =>  inp_feat(154), I1 =>  inp_feat(48), I2 =>  inp_feat(10), I3 =>  inp_feat(430), I4 =>  inp_feat(509), I5 =>  inp_feat(386), I6 =>  inp_feat(26), I7 =>  inp_feat(303)); 
C_37_S_2_L_0_inst : LUT8 generic map(INIT => "1111001111110101111000100000100011110011101010101000000010101010111101111111011100000000010000001111011110101010000000001010101000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_2_L_0_out, I0 =>  inp_feat(286), I1 =>  inp_feat(154), I2 =>  inp_feat(52), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_37_S_2_L_1_inst : LUT8 generic map(INIT => "1111000011110000101000001111010010110000100000001011000010000000111000001100000000000000101000001011000010000000101000000000000000000000101100000000000010000001000000001000000010000000100000000000000010010000000000001000000000000000000000001000000010000000") port map( O =>C_37_S_2_L_1_out, I0 =>  inp_feat(484), I1 =>  inp_feat(301), I2 =>  inp_feat(257), I3 =>  inp_feat(178), I4 =>  inp_feat(364), I5 =>  inp_feat(62), I6 =>  inp_feat(373), I7 =>  inp_feat(430)); 
C_37_S_2_L_2_inst : LUT8 generic map(INIT => "1111101011000000000000100000000011010101000000000000001000000000110010100100000011001010010000001100000000000000010000000100000011110111000000001000000000000000110101010000000000100000000000001010000010000000101000000000000000000000000000000000000000000000") port map( O =>C_37_S_2_L_2_out, I0 =>  inp_feat(39), I1 =>  inp_feat(399), I2 =>  inp_feat(150), I3 =>  inp_feat(310), I4 =>  inp_feat(273), I5 =>  inp_feat(157), I6 =>  inp_feat(316), I7 =>  inp_feat(280)); 
C_37_S_2_L_3_inst : LUT8 generic map(INIT => "1100010111001101101110110000000011001100010010010010000000000000010101011100010101110101010001000000010001000100010101010100010011000000110000001110000000000000110000001100000000000000000000001100000101000000011100000000000000000000000000000111000000000000") port map( O =>C_37_S_2_L_3_out, I0 =>  inp_feat(178), I1 =>  inp_feat(142), I2 =>  inp_feat(509), I3 =>  inp_feat(37), I4 =>  inp_feat(114), I5 =>  inp_feat(303), I6 =>  inp_feat(169), I7 =>  inp_feat(385)); 
C_37_S_2_L_4_inst : LUT8 generic map(INIT => "1111111111100000101000000000001011000100100000001100100000000000110011000000010011001100000000001100000000000000000010000000000011101010101010101000110010000000111100000000100011001100000001001000110000000000110010000000000010001000000000001000100000000000") port map( O =>C_37_S_2_L_4_out, I0 =>  inp_feat(301), I1 =>  inp_feat(307), I2 =>  inp_feat(74), I3 =>  inp_feat(77), I4 =>  inp_feat(382), I5 =>  inp_feat(367), I6 =>  inp_feat(169), I7 =>  inp_feat(286)); 
C_37_S_2_L_5_inst : LUT8 generic map(INIT => "1111111011000000110111000000000011111111100000001110110000000000111111000000000011110000000000000000000000000000000000000000000011001100100000001101000000000000100010001100000010001011010000001111110000000000111100000000000010101100000000000000000000000000") port map( O =>C_37_S_2_L_5_out, I0 =>  inp_feat(509), I1 =>  inp_feat(469), I2 =>  inp_feat(475), I3 =>  inp_feat(112), I4 =>  inp_feat(119), I5 =>  inp_feat(382), I6 =>  inp_feat(26), I7 =>  inp_feat(303)); 
C_37_S_2_L_6_inst : LUT8 generic map(INIT => "1011111111111000111110101111000000100010110000001101000011000000101010100000000011111011000000000010001000000000000000000000000011001010000000000000000000000000000000000000000000000000000000001100101100000000100010100000000000001010000000000000000000000000") port map( O =>C_37_S_2_L_6_out, I0 =>  inp_feat(364), I1 =>  inp_feat(56), I2 =>  inp_feat(29), I3 =>  inp_feat(216), I4 =>  inp_feat(31), I5 =>  inp_feat(430), I6 =>  inp_feat(119), I7 =>  inp_feat(470)); 
C_37_S_2_L_7_inst : LUT8 generic map(INIT => "1110111111001100110010001000110011101000110000001000000011000000101011001100111010100000100010001010000011001000000000001100100011100000110100000000000010000000000000001100000010000000010000001011000011100000101000001100000010110000111110000000000011001000") port map( O =>C_37_S_2_L_7_out, I0 =>  inp_feat(218), I1 =>  inp_feat(142), I2 =>  inp_feat(357), I3 =>  inp_feat(26), I4 =>  inp_feat(303), I5 =>  inp_feat(509), I6 =>  inp_feat(154), I7 =>  inp_feat(52)); 
C_37_S_3_L_0_inst : LUT8 generic map(INIT => "1111001111110101111000100000100011110011101010101000000010101010111101111111011100000000010000001111011110101010000000001010101000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_3_L_0_out, I0 =>  inp_feat(286), I1 =>  inp_feat(154), I2 =>  inp_feat(52), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_37_S_3_L_1_inst : LUT8 generic map(INIT => "1111110111110000111000001010000011110000100000001000000000000000010110001000000010001000101010001111100010000000100010000000000011011110110000001010000010000000100010001000100010100000000000001000110001000000100000001100000010001000100000001000000000000000") port map( O =>C_37_S_3_L_1_out, I0 =>  inp_feat(344), I1 =>  inp_feat(319), I2 =>  inp_feat(310), I3 =>  inp_feat(509), I4 =>  inp_feat(119), I5 =>  inp_feat(62), I6 =>  inp_feat(365), I7 =>  inp_feat(31)); 
C_37_S_3_L_2_inst : LUT8 generic map(INIT => "1111111010101000111011001000000011111100100100001110000110000000101100111011000011110000100000001011001010110000110000100000000010100010001000001010000010100000101000111011000110100000101000000010000000100000000000000000000000100000001100000000000000000000") port map( O =>C_37_S_3_L_2_out, I0 =>  inp_feat(48), I1 =>  inp_feat(509), I2 =>  inp_feat(142), I3 =>  inp_feat(303), I4 =>  inp_feat(216), I5 =>  inp_feat(151), I6 =>  inp_feat(253), I7 =>  inp_feat(430)); 
C_37_S_3_L_3_inst : LUT8 generic map(INIT => "1011100011101010000010001100100011010000000100001100000000000000111010101010001000000000000000001000000000000000000000000000000011001010100010101100000000000000100000000000000011000000000000001010101010000010100000000000000000000000000000000000000000000000") port map( O =>C_37_S_3_L_3_out, I0 =>  inp_feat(301), I1 =>  inp_feat(321), I2 =>  inp_feat(127), I3 =>  inp_feat(215), I4 =>  inp_feat(435), I5 =>  inp_feat(115), I6 =>  inp_feat(253), I7 =>  inp_feat(120)); 
C_37_S_3_L_4_inst : LUT8 generic map(INIT => "1110110011001100111001101010110010101010110000001010100010000000111011001100110010001001100011000000000000000000000000000000000011100000000000001010000010100000001000000000000010100000101000001100110001000100000001000000000000000000000000000000000000000000") port map( O =>C_37_S_3_L_4_out, I0 =>  inp_feat(247), I1 =>  inp_feat(222), I2 =>  inp_feat(273), I3 =>  inp_feat(203), I4 =>  inp_feat(301), I5 =>  inp_feat(372), I6 =>  inp_feat(399), I7 =>  inp_feat(6)); 
C_37_S_3_L_5_inst : LUT8 generic map(INIT => "1111111010001000110001000100010010001100100010000000110000000100110110000000100011010000010000001111100000000000000000000000000010001000000010000000000000000000100110000000000011110100000001000011000000000000000100000000000011110000000000001111000000000000") port map( O =>C_37_S_3_L_5_out, I0 =>  inp_feat(20), I1 =>  inp_feat(276), I2 =>  inp_feat(216), I3 =>  inp_feat(310), I4 =>  inp_feat(367), I5 =>  inp_feat(103), I6 =>  inp_feat(75), I7 =>  inp_feat(157)); 
C_37_S_3_L_6_inst : LUT8 generic map(INIT => "1111111011001000111111101010110111111000000010001000110010001100100100001000000010000000000000001011000000000000000000000000000010001000000000000000000000000000001110000000000000000000000000001001000000000000000000000000000011010000000000000000000000000000") port map( O =>C_37_S_3_L_6_out, I0 =>  inp_feat(161), I1 =>  inp_feat(218), I2 =>  inp_feat(5), I3 =>  inp_feat(142), I4 =>  inp_feat(108), I5 =>  inp_feat(328), I6 =>  inp_feat(358), I7 =>  inp_feat(57)); 
C_37_S_3_L_7_inst : LUT8 generic map(INIT => "1011110100000000001010000000000010101000100010001000100000000000111011000000000010101000000000001010100000000000101010000000000011001100110001001100110011000100100010001000100010001000100000000000000000000000000010000000000000000000000000000000100000000000") port map( O =>C_37_S_3_L_7_out, I0 =>  inp_feat(19), I1 =>  inp_feat(462), I2 =>  inp_feat(328), I3 =>  inp_feat(227), I4 =>  inp_feat(161), I5 =>  inp_feat(270), I6 =>  inp_feat(240), I7 =>  inp_feat(314)); 
C_37_S_4_L_0_inst : LUT8 generic map(INIT => "1111001111110101111000100000100011110011101010101000000010101010111101111111011100000000010000001111011110101010000000001010101000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_4_L_0_out, I0 =>  inp_feat(286), I1 =>  inp_feat(154), I2 =>  inp_feat(52), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_37_S_4_L_1_inst : LUT8 generic map(INIT => "1111110111110000111000001010000011110000100000001000000000000000010110001000000010001000101010001111100010000000100010000000000011011110110000001010000010000000100010001000100010100000000000001000110001000000100000001100000010001000100000001000000000000000") port map( O =>C_37_S_4_L_1_out, I0 =>  inp_feat(344), I1 =>  inp_feat(319), I2 =>  inp_feat(310), I3 =>  inp_feat(509), I4 =>  inp_feat(119), I5 =>  inp_feat(62), I6 =>  inp_feat(365), I7 =>  inp_feat(31)); 
C_37_S_4_L_2_inst : LUT8 generic map(INIT => "1011101110111010111110111000000010101010100010001010001000000000111000000000000011100010110000001010000000000000001000100000000000100110000000001100000000000000100010100000000010000000000000001000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_37_S_4_L_2_out, I0 =>  inp_feat(161), I1 =>  inp_feat(9), I2 =>  inp_feat(239), I3 =>  inp_feat(83), I4 =>  inp_feat(216), I5 =>  inp_feat(151), I6 =>  inp_feat(253), I7 =>  inp_feat(430)); 
C_37_S_4_L_3_inst : LUT8 generic map(INIT => "1111100010001110111100000100000000100010100000001110100010101010110010001000100011000000100000001100000010001000110000001000000011110010000000001111001000100010111010100000000010101010101000100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_4_L_3_out, I0 =>  inp_feat(218), I1 =>  inp_feat(50), I2 =>  inp_feat(475), I3 =>  inp_feat(383), I4 =>  inp_feat(26), I5 =>  inp_feat(303), I6 =>  inp_feat(485), I7 =>  inp_feat(240)); 
C_37_S_4_L_4_inst : LUT8 generic map(INIT => "1110100011111000111011101000000010100000101000100010001010100010111011101010101010101000000000100010000000100000100000000000001011101000101100111110110000000000101000100010001000101010001000001000100000000010000000100000000000000000000000100000100000000000") port map( O =>C_37_S_4_L_4_out, I0 =>  inp_feat(48), I1 =>  inp_feat(314), I2 =>  inp_feat(301), I3 =>  inp_feat(475), I4 =>  inp_feat(351), I5 =>  inp_feat(382), I6 =>  inp_feat(448), I7 =>  inp_feat(222)); 
C_37_S_4_L_5_inst : LUT8 generic map(INIT => "1110111000101000111010001100000010001010000000001110100011000000111011101010000000000000000000000010001000000000000000000000000000101000011000001000000011000000100000000000000010000000110000001111100011100000000000000000000000000000000000000000000000000000") port map( O =>C_37_S_4_L_5_out, I0 =>  inp_feat(301), I1 =>  inp_feat(303), I2 =>  inp_feat(50), I3 =>  inp_feat(455), I4 =>  inp_feat(347), I5 =>  inp_feat(382), I6 =>  inp_feat(26), I7 =>  inp_feat(245)); 
C_37_S_4_L_6_inst : LUT8 generic map(INIT => "1111010110100000110101000000000010100000101000000000000000000000110001001000000010000100100000001000110010000000000010000000000011111101110000000000010000000000110000000100000000000000000000001010110000000000000011000000000000001100000000000000100000000000") port map( O =>C_37_S_4_L_6_out, I0 =>  inp_feat(270), I1 =>  inp_feat(398), I2 =>  inp_feat(273), I3 =>  inp_feat(303), I4 =>  inp_feat(301), I5 =>  inp_feat(37), I6 =>  inp_feat(245), I7 =>  inp_feat(431)); 
C_37_S_4_L_7_inst : LUT8 generic map(INIT => "1110001011011110100000000000110011000000110000001100100011000000100000000100010010000000100000001000000011000000100000000000000010100000110000000000001010000000100000001100000000000000000000001010000011000010001000001100000011000000110000001100000000000000") port map( O =>C_37_S_4_L_7_out, I0 =>  inp_feat(303), I1 =>  inp_feat(301), I2 =>  inp_feat(142), I3 =>  inp_feat(494), I4 =>  inp_feat(207), I5 =>  inp_feat(379), I6 =>  inp_feat(77), I7 =>  inp_feat(203)); 
C_38_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000000000000000000010111010100000100000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000001000000000000000101010100000000000000000000000000000000000000000") port map( O =>C_38_S_0_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(316), I2 =>  inp_feat(470), I3 =>  inp_feat(371), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_38_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000001000000000000000000000001000001100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001110100110000001100000000000011110000000000000000000000000000000000000000000000000000000000000010") port map( O =>C_38_S_0_L_1_out, I0 =>  inp_feat(466), I1 =>  inp_feat(218), I2 =>  inp_feat(382), I3 =>  inp_feat(303), I4 =>  inp_feat(413), I5 =>  inp_feat(509), I6 =>  inp_feat(154), I7 =>  inp_feat(52)); 
C_38_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000100000000000000000011000001010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000100001000010000100010000110001010101110000000000000000000000000000000000000000110010000011000000110101") port map( O =>C_38_S_0_L_2_out, I0 =>  inp_feat(171), I1 =>  inp_feat(303), I2 =>  inp_feat(475), I3 =>  inp_feat(218), I4 =>  inp_feat(382), I5 =>  inp_feat(48), I6 =>  inp_feat(466), I7 =>  inp_feat(77)); 
C_38_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000100000000000000000011000001010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000100001000010000100010000110001010101110000000000000000000000000000000000000000110010000011000000110101") port map( O =>C_38_S_0_L_3_out, I0 =>  inp_feat(171), I1 =>  inp_feat(303), I2 =>  inp_feat(475), I3 =>  inp_feat(218), I4 =>  inp_feat(382), I5 =>  inp_feat(48), I6 =>  inp_feat(466), I7 =>  inp_feat(77)); 
C_38_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000100000000000000000011000001010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000100001000010000100010000110001010101110000000000000000000000000000000000000000110010000011000000110101") port map( O =>C_38_S_0_L_4_out, I0 =>  inp_feat(171), I1 =>  inp_feat(303), I2 =>  inp_feat(475), I3 =>  inp_feat(218), I4 =>  inp_feat(382), I5 =>  inp_feat(48), I6 =>  inp_feat(466), I7 =>  inp_feat(77)); 
C_38_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000100000000000000000011000001010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000100001000010000100010000110001010101110000000000000000000000000000000000000000110010000011000000110101") port map( O =>C_38_S_0_L_5_out, I0 =>  inp_feat(171), I1 =>  inp_feat(303), I2 =>  inp_feat(475), I3 =>  inp_feat(218), I4 =>  inp_feat(382), I5 =>  inp_feat(48), I6 =>  inp_feat(466), I7 =>  inp_feat(77)); 
C_38_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000100000000000000000011000001010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000100001000010000100010000110001010101110000000000000000000000000000000000000000110010000011000000110101") port map( O =>C_38_S_0_L_6_out, I0 =>  inp_feat(171), I1 =>  inp_feat(303), I2 =>  inp_feat(475), I3 =>  inp_feat(218), I4 =>  inp_feat(382), I5 =>  inp_feat(48), I6 =>  inp_feat(466), I7 =>  inp_feat(77)); 
C_38_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000100000000000000000011000001010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000100001000010000100010000110001010101110000000000000000000000000000000000000000110010000011000000110101") port map( O =>C_38_S_0_L_7_out, I0 =>  inp_feat(171), I1 =>  inp_feat(303), I2 =>  inp_feat(475), I3 =>  inp_feat(218), I4 =>  inp_feat(382), I5 =>  inp_feat(48), I6 =>  inp_feat(466), I7 =>  inp_feat(77)); 
C_38_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000000000000000000010111010100000100000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000001000000000000000101010100000000000000000000000000000000000000000") port map( O =>C_38_S_1_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(316), I2 =>  inp_feat(470), I3 =>  inp_feat(371), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_38_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000001000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000000000010000000100010001010101010001000100000000000000000000000000000000000000000000000000010001000000000") port map( O =>C_38_S_1_L_1_out, I0 =>  inp_feat(286), I1 =>  inp_feat(218), I2 =>  inp_feat(201), I3 =>  inp_feat(136), I4 =>  inp_feat(303), I5 =>  inp_feat(142), I6 =>  inp_feat(154), I7 =>  inp_feat(52)); 
C_38_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000100000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000101000010000100110001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_1_L_2_out, I0 =>  inp_feat(382), I1 =>  inp_feat(286), I2 =>  inp_feat(41), I3 =>  inp_feat(218), I4 =>  inp_feat(509), I5 =>  inp_feat(420), I6 =>  inp_feat(9), I7 =>  inp_feat(307)); 
C_38_S_1_L_3_inst : LUT8 generic map(INIT => "0000000100000111000000000000001000000010000000011010001000000011000000010000000000000000000000000000000000000000000000000000000000010001000101110000000000000010000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_1_L_3_out, I0 =>  inp_feat(303), I1 =>  inp_feat(218), I2 =>  inp_feat(142), I3 =>  inp_feat(225), I4 =>  inp_feat(425), I5 =>  inp_feat(474), I6 =>  inp_feat(178), I7 =>  inp_feat(37)); 
C_38_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000001000000010000000000000000000000000000000000001010000000000010000100000000000000010000000000000000010000000000000000000000000000010000000000000011000000000000001100000000000011110000000000000000000100010001000101010000000100010001000000010001") port map( O =>C_38_S_1_L_4_out, I0 =>  inp_feat(222), I1 =>  inp_feat(218), I2 =>  inp_feat(247), I3 =>  inp_feat(303), I4 =>  inp_feat(212), I5 =>  inp_feat(98), I6 =>  inp_feat(78), I7 =>  inp_feat(77)); 
C_38_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000001100000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000101000011110000000000101111000000010000000000000000000000000000000000100000000000000000000000000000") port map( O =>C_38_S_1_L_5_out, I0 =>  inp_feat(61), I1 =>  inp_feat(218), I2 =>  inp_feat(48), I3 =>  inp_feat(425), I4 =>  inp_feat(494), I5 =>  inp_feat(382), I6 =>  inp_feat(180), I7 =>  inp_feat(52)); 
C_38_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000100000100000000000001010001100000010000000000000001010100000000000100000000000000010101000000000001000100000000000000000000000000000000000000000001000100011000000100000000000000010001000100000000000100000000000100010000000000010000000000000") port map( O =>C_38_S_1_L_6_out, I0 =>  inp_feat(160), I1 =>  inp_feat(142), I2 =>  inp_feat(323), I3 =>  inp_feat(82), I4 =>  inp_feat(13), I5 =>  inp_feat(407), I6 =>  inp_feat(358), I7 =>  inp_feat(370)); 
C_38_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000000000000000000010000000000000001100000100000000100001000000100000000000100010001100100000000000010000000000000001001000000000000000000000001000000000000000000011000000010000001000000000000000110000001000000011000000") port map( O =>C_38_S_1_L_7_out, I0 =>  inp_feat(177), I1 =>  inp_feat(388), I2 =>  inp_feat(5), I3 =>  inp_feat(239), I4 =>  inp_feat(227), I5 =>  inp_feat(323), I6 =>  inp_feat(303), I7 =>  inp_feat(236)); 
C_38_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000000000000000000010111010100000100000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000001000000000000000101010100000000000000000000000000000000000000000") port map( O =>C_38_S_2_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(316), I2 =>  inp_feat(470), I3 =>  inp_feat(371), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_38_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000001000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000000000010000000100010001010101010001000100000000000000000000000000000000000000000000000000010001000000000") port map( O =>C_38_S_2_L_1_out, I0 =>  inp_feat(286), I1 =>  inp_feat(218), I2 =>  inp_feat(201), I3 =>  inp_feat(136), I4 =>  inp_feat(303), I5 =>  inp_feat(142), I6 =>  inp_feat(154), I7 =>  inp_feat(52)); 
C_38_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000100000000000000000000100000110011101100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000100011111000110001100110011000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_2_L_2_out, I0 =>  inp_feat(475), I1 =>  inp_feat(112), I2 =>  inp_feat(473), I3 =>  inp_feat(218), I4 =>  inp_feat(364), I5 =>  inp_feat(420), I6 =>  inp_feat(9), I7 =>  inp_feat(307)); 
C_38_S_2_L_3_inst : LUT8 generic map(INIT => "1010001100000000000000000000000000010001000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_2_L_3_out, I0 =>  inp_feat(238), I1 =>  inp_feat(218), I2 =>  inp_feat(470), I3 =>  inp_feat(31), I4 =>  inp_feat(345), I5 =>  inp_feat(9), I6 =>  inp_feat(178), I7 =>  inp_feat(237)); 
C_38_S_2_L_4_inst : LUT8 generic map(INIT => "0000000001010011000000000000000000000000000000010000000000000000000000000000001100000000000000000000000010010001000000000000000100000000000001110000000000000000000000000000000100000000000000010001000100000011000000000000000000000000000001010000000000000000") port map( O =>C_38_S_2_L_4_out, I0 =>  inp_feat(218), I1 =>  inp_feat(448), I2 =>  inp_feat(245), I3 =>  inp_feat(509), I4 =>  inp_feat(17), I5 =>  inp_feat(134), I6 =>  inp_feat(307), I7 =>  inp_feat(37)); 
C_38_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000010000001000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000100010000001100110011001100000000000000000000000000000000000100000000000000010000000000000000000000000000001000000000000000") port map( O =>C_38_S_2_L_5_out, I0 =>  inp_feat(218), I1 =>  inp_feat(68), I2 =>  inp_feat(342), I3 =>  inp_feat(174), I4 =>  inp_feat(386), I5 =>  inp_feat(270), I6 =>  inp_feat(64), I7 =>  inp_feat(77)); 
C_38_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000010001000000000000000000000000000000010000000000010000000100010001000100000000000101000000000100000000000000000011000100000000000100000000000000") port map( O =>C_38_S_2_L_6_out, I0 =>  inp_feat(218), I1 =>  inp_feat(237), I2 =>  inp_feat(200), I3 =>  inp_feat(446), I4 =>  inp_feat(452), I5 =>  inp_feat(448), I6 =>  inp_feat(227), I7 =>  inp_feat(382)); 
C_38_S_2_L_7_inst : LUT8 generic map(INIT => "0010000000011100000000000000000000000000000010000000000000000000000010001000100000000000000000000100000000001000000000000000000000000000011100100000000000000000010000000000000000000000000000000000000000001000010000000000000001000000100000000000000000000000") port map( O =>C_38_S_2_L_7_out, I0 =>  inp_feat(162), I1 =>  inp_feat(112), I2 =>  inp_feat(37), I3 =>  inp_feat(77), I4 =>  inp_feat(178), I5 =>  inp_feat(470), I6 =>  inp_feat(480), I7 =>  inp_feat(344)); 
C_38_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000000000000000000010111010100000100000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000001000000000000000101010100000000000000000000000000000000000000000") port map( O =>C_38_S_3_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(316), I2 =>  inp_feat(470), I3 =>  inp_feat(371), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_38_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000001000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000000000010000000100010001010101010001000100000000000000000000000000000000000000000000000000010001000000000") port map( O =>C_38_S_3_L_1_out, I0 =>  inp_feat(286), I1 =>  inp_feat(218), I2 =>  inp_feat(201), I3 =>  inp_feat(136), I4 =>  inp_feat(303), I5 =>  inp_feat(142), I6 =>  inp_feat(154), I7 =>  inp_feat(52)); 
C_38_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000001000100010101100000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000101010101000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_3_L_2_out, I0 =>  inp_feat(160), I1 =>  inp_feat(469), I2 =>  inp_feat(41), I3 =>  inp_feat(329), I4 =>  inp_feat(420), I5 =>  inp_feat(26), I6 =>  inp_feat(9), I7 =>  inp_feat(372)); 
C_38_S_3_L_3_inst : LUT8 generic map(INIT => "0100011100000000000001010000000000000100000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_3_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(228), I2 =>  inp_feat(218), I3 =>  inp_feat(508), I4 =>  inp_feat(470), I5 =>  inp_feat(9), I6 =>  inp_feat(178), I7 =>  inp_feat(359)); 
C_38_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000010000000101001101000000100000011100000001000001110000000000000001000001110000100100000010010000010000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000") port map( O =>C_38_S_3_L_4_out, I0 =>  inp_feat(303), I1 =>  inp_feat(7), I2 =>  inp_feat(295), I3 =>  inp_feat(434), I4 =>  inp_feat(301), I5 =>  inp_feat(333), I6 =>  inp_feat(87), I7 =>  inp_feat(287)); 
C_38_S_3_L_5_inst : LUT8 generic map(INIT => "0000001000000000000000000000000000000000000001000000001100000000000000000000000000000000000000000000000000000000000000000000000001000111000000001001000000000000000101110000000000100001000000000000000000000000000000000000000001000000000000000000000000000000") port map( O =>C_38_S_3_L_5_out, I0 =>  inp_feat(48), I1 =>  inp_feat(469), I2 =>  inp_feat(448), I3 =>  inp_feat(284), I4 =>  inp_feat(5), I5 =>  inp_feat(77), I6 =>  inp_feat(270), I7 =>  inp_feat(435)); 
C_38_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000011010000100001000000000000000000100011000000000000000000000000000000110000000000000000000000100010001000000000000000000000000000001100000010100000000000000010000011000000111100000000000000000000000000000000000000000000101000000000000011100000") port map( O =>C_38_S_3_L_6_out, I0 =>  inp_feat(5), I1 =>  inp_feat(239), I2 =>  inp_feat(425), I3 =>  inp_feat(298), I4 =>  inp_feat(108), I5 =>  inp_feat(414), I6 =>  inp_feat(370), I7 =>  inp_feat(358)); 
C_38_S_3_L_7_inst : LUT8 generic map(INIT => "0000000100000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010011111100000101000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_38_S_3_L_7_out, I0 =>  inp_feat(509), I1 =>  inp_feat(372), I2 =>  inp_feat(52), I3 =>  inp_feat(465), I4 =>  inp_feat(247), I5 =>  inp_feat(286), I6 =>  inp_feat(178), I7 =>  inp_feat(218)); 
C_38_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000000000000000000010111010100000100000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000001000000000000000101010100000000000000000000000000000000000000000") port map( O =>C_38_S_4_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(316), I2 =>  inp_feat(470), I3 =>  inp_feat(371), I4 =>  inp_feat(218), I5 =>  inp_feat(178), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_38_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000100110101000000010001000000010001000100000001000000000001010100000001010") port map( O =>C_38_S_4_L_1_out, I0 =>  inp_feat(388), I1 =>  inp_feat(451), I2 =>  inp_feat(414), I3 =>  inp_feat(310), I4 =>  inp_feat(303), I5 =>  inp_feat(364), I6 =>  inp_feat(48), I7 =>  inp_feat(52)); 
C_38_S_4_L_2_inst : LUT8 generic map(INIT => "0000001100000001001100110000000001000111000000000011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000") port map( O =>C_38_S_4_L_2_out, I0 =>  inp_feat(222), I1 =>  inp_feat(303), I2 =>  inp_feat(218), I3 =>  inp_feat(351), I4 =>  inp_feat(257), I5 =>  inp_feat(457), I6 =>  inp_feat(120), I7 =>  inp_feat(12)); 
C_38_S_4_L_3_inst : LUT8 generic map(INIT => "0000000001000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000001000100110100010000000001000001010000001100000000000000000000000000000011010000000000000000000000000000010000000000000000000000") port map( O =>C_38_S_4_L_3_out, I0 =>  inp_feat(509), I1 =>  inp_feat(419), I2 =>  inp_feat(156), I3 =>  inp_feat(218), I4 =>  inp_feat(58), I5 =>  inp_feat(466), I6 =>  inp_feat(484), I7 =>  inp_feat(161)); 
C_38_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000001110000000000000000000000000000000000000100000000100000000000000001000000000010001000000000000000010000000000000100000000000000011100000000010001010000000001000101000000000000000000000000000000010000000000010000000000000000010100000000") port map( O =>C_38_S_4_L_4_out, I0 =>  inp_feat(382), I1 =>  inp_feat(157), I2 =>  inp_feat(77), I3 =>  inp_feat(215), I4 =>  inp_feat(53), I5 =>  inp_feat(212), I6 =>  inp_feat(13), I7 =>  inp_feat(358)); 
C_38_S_4_L_5_inst : LUT8 generic map(INIT => "0001000000000001000000000000000000000000000000010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010000010100000011010101000000000000010011000000111101010000000000000000000000000000000000000000100011000000000001000000") port map( O =>C_38_S_4_L_5_out, I0 =>  inp_feat(72), I1 =>  inp_feat(328), I2 =>  inp_feat(398), I3 =>  inp_feat(161), I4 =>  inp_feat(171), I5 =>  inp_feat(11), I6 =>  inp_feat(95), I7 =>  inp_feat(218)); 
C_38_S_4_L_6_inst : LUT8 generic map(INIT => "0000001000001010000000000000000010001010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000101011000010110000000000000000000010100000101000000000000000000000000000000000000000010000000000000000000000000000000000000000") port map( O =>C_38_S_4_L_6_out, I0 =>  inp_feat(275), I1 =>  inp_feat(469), I2 =>  inp_feat(420), I3 =>  inp_feat(466), I4 =>  inp_feat(109), I5 =>  inp_feat(174), I6 =>  inp_feat(287), I7 =>  inp_feat(310)); 
C_38_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000100000100000000000000000000000000000000000000000000001000000000100000000000000000000010000000001000000000000010000000100000001010000011000100000000001100000010100000100000001000000010000000") port map( O =>C_38_S_4_L_7_out, I0 =>  inp_feat(200), I1 =>  inp_feat(112), I2 =>  inp_feat(314), I3 =>  inp_feat(468), I4 =>  inp_feat(373), I5 =>  inp_feat(358), I6 =>  inp_feat(239), I7 =>  inp_feat(448)); 
C_39_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000000000000000000000000100000000000101010000000100000000000000000000010000000000000000000000000000010001000000000000000000000000000000000000000000000100000000000001010100000000000000000000000000000000000000000") port map( O =>C_39_S_0_L_0_out, I0 =>  inp_feat(315), I1 =>  inp_feat(204), I2 =>  inp_feat(48), I3 =>  inp_feat(103), I4 =>  inp_feat(218), I5 =>  inp_feat(249), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_39_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000010000000001100000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000001000100010101000000100001111000000001000100000000000100010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_0_L_1_out, I0 =>  inp_feat(12), I1 =>  inp_feat(394), I2 =>  inp_feat(509), I3 =>  inp_feat(161), I4 =>  inp_feat(86), I5 =>  inp_feat(196), I6 =>  inp_feat(62), I7 =>  inp_feat(365)); 
C_39_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000011000000000000000100010001000000000000000000000000000000010000000100110000000000000000000100000101000000000000000000000001000000010000000000000001000000") port map( O =>C_39_S_0_L_2_out, I0 =>  inp_feat(365), I1 =>  inp_feat(26), I2 =>  inp_feat(180), I3 =>  inp_feat(509), I4 =>  inp_feat(451), I5 =>  inp_feat(303), I6 =>  inp_feat(142), I7 =>  inp_feat(430)); 
C_39_S_0_L_3_inst : LUT8 generic map(INIT => "0000000001001010001000000001010000000000100000000000101010001111000000000000000000000000000000000000000000000000000000000000010010000000110010000000000000001111000000000000110100000000000011110000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_0_L_3_out, I0 =>  inp_feat(81), I1 =>  inp_feat(189), I2 =>  inp_feat(382), I3 =>  inp_feat(142), I4 =>  inp_feat(303), I5 =>  inp_feat(247), I6 =>  inp_feat(314), I7 =>  inp_feat(227)); 
C_39_S_0_L_4_inst : LUT8 generic map(INIT => "0000000010000000001000000010000000000000100000000010000000000000101000001010000000100000001000100000000000000000000100100000000000001010101000000000000010100000000000001000000000000000100000001000000010100000000000000000000010000000000000000000000000000000") port map( O =>C_39_S_0_L_4_out, I0 =>  inp_feat(388), I1 =>  inp_feat(88), I2 =>  inp_feat(331), I3 =>  inp_feat(430), I4 =>  inp_feat(344), I5 =>  inp_feat(180), I6 =>  inp_feat(247), I7 =>  inp_feat(455)); 
C_39_S_0_L_5_inst : LUT8 generic map(INIT => "0000010000001101000001010001110100000000000011000000101000001100000000001100110000000000000011010100100001001110000000000000110000000000000000000000000000001000000000000000100000000000000000000100000011100100000000000000000000000000000000000000000000000000") port map( O =>C_39_S_0_L_5_out, I0 =>  inp_feat(229), I1 =>  inp_feat(5), I2 =>  inp_feat(386), I3 =>  inp_feat(382), I4 =>  inp_feat(333), I5 =>  inp_feat(40), I6 =>  inp_feat(301), I7 =>  inp_feat(470)); 
C_39_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000110000011000000000000000000000000000000000000000000000000000000001000000000000010010001000000000001000000000100000000000101000001010000110100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_0_L_6_out, I0 =>  inp_feat(77), I1 =>  inp_feat(430), I2 =>  inp_feat(287), I3 =>  inp_feat(40), I4 =>  inp_feat(386), I5 =>  inp_feat(298), I6 =>  inp_feat(26), I7 =>  inp_feat(218)); 
C_39_S_0_L_7_inst : LUT8 generic map(INIT => "0001000100000000110100000000000001010110000000000111000101010010010100000000000010010000000000000001000000000000100000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_0_L_7_out, I0 =>  inp_feat(142), I1 =>  inp_feat(469), I2 =>  inp_feat(145), I3 =>  inp_feat(25), I4 =>  inp_feat(48), I5 =>  inp_feat(77), I6 =>  inp_feat(354), I7 =>  inp_feat(286)); 
C_39_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000000000000000000000000100000000000101010000000100000000000000000000010000000000000000000000000000010001000000000000000000000000000000000000000000000100000000000001010100000000000000000000000000000000000000000") port map( O =>C_39_S_1_L_0_out, I0 =>  inp_feat(315), I1 =>  inp_feat(204), I2 =>  inp_feat(48), I3 =>  inp_feat(103), I4 =>  inp_feat(218), I5 =>  inp_feat(249), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_39_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000010000000001100000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000001000100010101000000100001111000000000000000000000000000000000000000010001000000000001000100000000000000000000000000000000000") port map( O =>C_39_S_1_L_1_out, I0 =>  inp_feat(12), I1 =>  inp_feat(394), I2 =>  inp_feat(509), I3 =>  inp_feat(161), I4 =>  inp_feat(86), I5 =>  inp_feat(62), I6 =>  inp_feat(196), I7 =>  inp_feat(365)); 
C_39_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000001011100000000000001000000000000010010000000000001110010000000000101000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000") port map( O =>C_39_S_1_L_2_out, I0 =>  inp_feat(249), I1 =>  inp_feat(298), I2 =>  inp_feat(279), I3 =>  inp_feat(131), I4 =>  inp_feat(413), I5 =>  inp_feat(509), I6 =>  inp_feat(430), I7 =>  inp_feat(286)); 
C_39_S_1_L_3_inst : LUT8 generic map(INIT => "0001000100000000000000000000000001000101000010010000000000000000100100010000000000000000000000000001010111110111000011000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_1_L_3_out, I0 =>  inp_feat(218), I1 =>  inp_feat(15), I2 =>  inp_feat(301), I3 =>  inp_feat(105), I4 =>  inp_feat(56), I5 =>  inp_feat(382), I6 =>  inp_feat(303), I7 =>  inp_feat(26)); 
C_39_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000001000001000010110001100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000010000010101001000000000000000000000000000000010000000000110000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_1_L_4_out, I0 =>  inp_feat(220), I1 =>  inp_feat(273), I2 =>  inp_feat(301), I3 =>  inp_feat(34), I4 =>  inp_feat(386), I5 =>  inp_feat(26), I6 =>  inp_feat(429), I7 =>  inp_feat(364)); 
C_39_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000010000000000000000000001110000001100000000000000000000001100000111000000000000000000000100110000000000000000000000000000000001000100000001000000010000001110000011000000000000000000000000000000100000000000000000000000000000001000100000000000000000") port map( O =>C_39_S_1_L_5_out, I0 =>  inp_feat(307), I1 =>  inp_feat(509), I2 =>  inp_feat(109), I3 =>  inp_feat(302), I4 =>  inp_feat(216), I5 =>  inp_feat(247), I6 =>  inp_feat(344), I7 =>  inp_feat(475)); 
C_39_S_1_L_6_inst : LUT8 generic map(INIT => "0000000100000000000100011101000100000100101100100101000001000000000000000000000100000000010100010100000010110100010100001111010100000000000000000000000000100000000001001000000000000000000000000000000000000000000000000000000000000000001100000000000000100000") port map( O =>C_39_S_1_L_6_out, I0 =>  inp_feat(77), I1 =>  inp_feat(469), I2 =>  inp_feat(198), I3 =>  inp_feat(19), I4 =>  inp_feat(386), I5 =>  inp_feat(301), I6 =>  inp_feat(334), I7 =>  inp_feat(351)); 
C_39_S_1_L_7_inst : LUT8 generic map(INIT => "0001000000000010000000001101010000000000000000001001100011010000000000000000001000000000010100000000000000000000010100000001000000000000010000000000000001010000000000000100000010011100110100000000000001000000000000000100000000000000110000000101100011010000") port map( O =>C_39_S_1_L_7_out, I0 =>  inp_feat(77), I1 =>  inp_feat(430), I2 =>  inp_feat(371), I3 =>  inp_feat(386), I4 =>  inp_feat(52), I5 =>  inp_feat(301), I6 =>  inp_feat(221), I7 =>  inp_feat(334)); 
C_39_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000000000000000000000000100000000000101010000000100000000000000000000010000000000000000000000000000010001000000000000000000000000000000000000000000000100000000000001010100000000000000000000000000000000000000000") port map( O =>C_39_S_2_L_0_out, I0 =>  inp_feat(315), I1 =>  inp_feat(204), I2 =>  inp_feat(48), I3 =>  inp_feat(103), I4 =>  inp_feat(218), I5 =>  inp_feat(249), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_39_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000001000100010001010100010001000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000") port map( O =>C_39_S_2_L_1_out, I0 =>  inp_feat(151), I1 =>  inp_feat(26), I2 =>  inp_feat(244), I3 =>  inp_feat(497), I4 =>  inp_feat(382), I5 =>  inp_feat(62), I6 =>  inp_feat(196), I7 =>  inp_feat(365)); 
C_39_S_2_L_2_inst : LUT8 generic map(INIT => "1101001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_2_L_2_out, I0 =>  inp_feat(247), I1 =>  inp_feat(321), I2 =>  inp_feat(115), I3 =>  inp_feat(110), I4 =>  inp_feat(30), I5 =>  inp_feat(266), I6 =>  inp_feat(353), I7 =>  inp_feat(119)); 
C_39_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000001000000000000000000001101001010110001000000010011000000000000000000000000000000000000000000000001000000000001000000000010100100000000000000000000010000010011001100001000000000010000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_2_L_3_out, I0 =>  inp_feat(301), I1 =>  inp_feat(142), I2 =>  inp_feat(86), I3 =>  inp_feat(448), I4 =>  inp_feat(128), I5 =>  inp_feat(509), I6 =>  inp_feat(154), I7 =>  inp_feat(430)); 
C_39_S_2_L_4_inst : LUT8 generic map(INIT => "0001000000000000000000000000000001010100000000000100000000000000000011010000000000000000000000011111111100000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000100000000000001000000000100000101000000001000000000000000") port map( O =>C_39_S_2_L_4_out, I0 =>  inp_feat(53), I1 =>  inp_feat(480), I2 =>  inp_feat(301), I3 =>  inp_feat(56), I4 =>  inp_feat(371), I5 =>  inp_feat(386), I6 =>  inp_feat(142), I7 =>  inp_feat(419)); 
C_39_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000001000010100010000000000000000000000000000110000000000000010000001000011011001010100010000000000000000000001010000000000000111000000000000111100100010000011110000000010001111000000000000000110000000010100010001000100000001000000000000000100000000") port map( O =>C_39_S_2_L_5_out, I0 =>  inp_feat(53), I1 =>  inp_feat(301), I2 =>  inp_feat(19), I3 =>  inp_feat(156), I4 =>  inp_feat(218), I5 =>  inp_feat(217), I6 =>  inp_feat(475), I7 =>  inp_feat(212)); 
C_39_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000010111010000010000010000000000000100100000000000000010000000000000000000000000000000100000010000000000000000000001011100000111000100110100001100011000000000000000010000000100000000000000000000000000000000010000000000000000000000000000010000") port map( O =>C_39_S_2_L_6_out, I0 =>  inp_feat(301), I1 =>  inp_feat(90), I2 =>  inp_feat(386), I3 =>  inp_feat(444), I4 =>  inp_feat(222), I5 =>  inp_feat(344), I6 =>  inp_feat(180), I7 =>  inp_feat(247)); 
C_39_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000010000000000000011000000000000000100000000000000110000000000000000000000100000001100100100000001110000001000000011001000000000000100000000000000110010001000001000000000000000001100000000000000000000000000100000000001000000001110000000000000110000") port map( O =>C_39_S_2_L_7_out, I0 =>  inp_feat(57), I1 =>  inp_feat(340), I2 =>  inp_feat(145), I3 =>  inp_feat(303), I4 =>  inp_feat(41), I5 =>  inp_feat(494), I6 =>  inp_feat(211), I7 =>  inp_feat(290)); 
C_39_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000000000000000000000000100000000000101010000000100000000000000000000010000000000000000000000000000010001000000000000000000000000000000000000000000000100000000000001010100000000000000000000000000000000000000000") port map( O =>C_39_S_3_L_0_out, I0 =>  inp_feat(315), I1 =>  inp_feat(204), I2 =>  inp_feat(48), I3 =>  inp_feat(103), I4 =>  inp_feat(218), I5 =>  inp_feat(249), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_39_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000001000000000000000000010000000000000000000000000000000000100000010100000000000000000000111101011111000000000000000000000001000000000000000000000000000001000100010000000000000000000010001100000101001000100000000000001101100001010000000000000000") port map( O =>C_39_S_3_L_1_out, I0 =>  inp_feat(450), I1 =>  inp_feat(301), I2 =>  inp_feat(218), I3 =>  inp_feat(189), I4 =>  inp_feat(160), I5 =>  inp_feat(427), I6 =>  inp_feat(142), I7 =>  inp_feat(71)); 
C_39_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000010000000010000000000000001100000011000000010000000000000000000000000000000000000000000000010000000100000001000001000000000000001110000000110000000000000001100000010000010100000000000000000000000000000010000000000000000000000001000000000000") port map( O =>C_39_S_3_L_2_out, I0 =>  inp_feat(303), I1 =>  inp_feat(509), I2 =>  inp_feat(26), I3 =>  inp_feat(386), I4 =>  inp_feat(52), I5 =>  inp_feat(19), I6 =>  inp_feat(115), I7 =>  inp_feat(430)); 
C_39_S_3_L_3_inst : LUT8 generic map(INIT => "0000001000000000001000100000000000001010000000001010101000000000000000000000000000000000000000000000000000000000000010000000000010100000000000001010001000000000001000000000000010101010000000000000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_39_S_3_L_3_out, I0 =>  inp_feat(39), I1 =>  inp_feat(227), I2 =>  inp_feat(212), I3 =>  inp_feat(240), I4 =>  inp_feat(303), I5 =>  inp_feat(247), I6 =>  inp_feat(314), I7 =>  inp_feat(290)); 
C_39_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000101000000000000000000000000001000010000000000001001000000000000010000000000000000000000000000000000000000000010110000000001000111111000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_3_L_4_out, I0 =>  inp_feat(301), I1 =>  inp_feat(358), I2 =>  inp_feat(394), I3 =>  inp_feat(154), I4 =>  inp_feat(227), I5 =>  inp_feat(216), I6 =>  inp_feat(180), I7 =>  inp_feat(448)); 
C_39_S_3_L_5_inst : LUT8 generic map(INIT => "0000001000111010000000000000100000000000000000000000000000000000101110101010101010100000000010000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_3_L_5_out, I0 =>  inp_feat(238), I1 =>  inp_feat(19), I2 =>  inp_feat(473), I3 =>  inp_feat(204), I4 =>  inp_feat(262), I5 =>  inp_feat(131), I6 =>  inp_feat(430), I7 =>  inp_feat(154)); 
C_39_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000101010000000001010101000000100000111000001000010001010000000000000000000000000000010101100000000001000000010000000100000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_3_L_6_out, I0 =>  inp_feat(354), I1 =>  inp_feat(5), I2 =>  inp_feat(273), I3 =>  inp_feat(77), I4 =>  inp_feat(37), I5 =>  inp_feat(301), I6 =>  inp_feat(83), I7 =>  inp_feat(111)); 
C_39_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000010001000000001000000100000000000100010000000000000000000000000000110000001000000000010000000000010001000001000100010000000000000001000100000100000001010000010000000100000000000000000000000000000000000000000000000100000000000000010") port map( O =>C_39_S_3_L_7_out, I0 =>  inp_feat(151), I1 =>  inp_feat(48), I2 =>  inp_feat(161), I3 =>  inp_feat(218), I4 =>  inp_feat(229), I5 =>  inp_feat(386), I6 =>  inp_feat(13), I7 =>  inp_feat(413)); 
C_39_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000000000000000000000000100000000000101010000000100000000000000000000010000000000000000000000000000010001000000000000000000000000000000000000000000000100000000000001010100000000000000000000000000000000000000000") port map( O =>C_39_S_4_L_0_out, I0 =>  inp_feat(315), I1 =>  inp_feat(204), I2 =>  inp_feat(48), I3 =>  inp_feat(103), I4 =>  inp_feat(218), I5 =>  inp_feat(249), I6 =>  inp_feat(509), I7 =>  inp_feat(257)); 
C_39_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000001000000000001000100000000000000100100010000010001000000000011001100000000000100110000000000000000000000000000000000110000000000010000000000100000000000000000000000010010000100100010001000000011000000000000001100") port map( O =>C_39_S_4_L_1_out, I0 =>  inp_feat(227), I1 =>  inp_feat(151), I2 =>  inp_feat(399), I3 =>  inp_feat(43), I4 =>  inp_feat(307), I5 =>  inp_feat(364), I6 =>  inp_feat(77), I7 =>  inp_feat(71)); 
C_39_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000001000001000000000101000000000000000000000000000000000001100101000100010101010000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_4_L_2_out, I0 =>  inp_feat(26), I1 =>  inp_feat(382), I2 =>  inp_feat(112), I3 =>  inp_feat(271), I4 =>  inp_feat(161), I5 =>  inp_feat(286), I6 =>  inp_feat(430), I7 =>  inp_feat(240)); 
C_39_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000000000000000000000000000010000000000000000110000000010000000000000000000000000010000000000000000000000000000000000000000000000100000001000000000000100010100000001000111101000110000110000001011100011110000001100000111") port map( O =>C_39_S_4_L_3_out, I0 =>  inp_feat(98), I1 =>  inp_feat(247), I2 =>  inp_feat(358), I3 =>  inp_feat(430), I4 =>  inp_feat(413), I5 =>  inp_feat(121), I6 =>  inp_feat(509), I7 =>  inp_feat(218)); 
C_39_S_4_L_4_inst : LUT8 generic map(INIT => "0010100101110100011100000101010000010000000000000100000000000100000000000000000000000000000000001000000010000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_4_L_4_out, I0 =>  inp_feat(340), I1 =>  inp_feat(430), I2 =>  inp_feat(371), I3 =>  inp_feat(301), I4 =>  inp_feat(373), I5 =>  inp_feat(347), I6 =>  inp_feat(415), I7 =>  inp_feat(390)); 
C_39_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000001010000000000000000000101000000000001000100000001000000000000000000000000000000000000100100000000000100010000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000011110000000000000000000000000000") port map( O =>C_39_S_4_L_5_out, I0 =>  inp_feat(374), I1 =>  inp_feat(20), I2 =>  inp_feat(227), I3 =>  inp_feat(425), I4 =>  inp_feat(430), I5 =>  inp_feat(142), I6 =>  inp_feat(344), I7 =>  inp_feat(111)); 
C_39_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000100010000000100000000001010000101000010001000000000000000000000000000000000000000000010000000000000000000000010011000000000111001001010000001100010000000001110011000010010000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_4_L_6_out, I0 =>  inp_feat(469), I1 =>  inp_feat(142), I2 =>  inp_feat(475), I3 =>  inp_feat(34), I4 =>  inp_feat(450), I5 =>  inp_feat(386), I6 =>  inp_feat(26), I7 =>  inp_feat(303)); 
C_39_S_4_L_7_inst : LUT8 generic map(INIT => "0111010001010000010100001111100000000000000000000000000010000000010000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_39_S_4_L_7_out, I0 =>  inp_feat(142), I1 =>  inp_feat(303), I2 =>  inp_feat(151), I3 =>  inp_feat(204), I4 =>  inp_feat(57), I5 =>  inp_feat(103), I6 =>  inp_feat(351), I7 =>  inp_feat(119)); 
C_40_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000100000001000001010000000000000001000000000000010000000000000000000000010111010101000000000000010100000000010000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000") port map( O =>C_40_S_0_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(57), I2 =>  inp_feat(204), I3 =>  inp_feat(496), I4 =>  inp_feat(27), I5 =>  inp_feat(484), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_40_S_0_L_1_inst : LUT8 generic map(INIT => "0000000010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000110100000100000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_0_L_1_out, I0 =>  inp_feat(134), I1 =>  inp_feat(29), I2 =>  inp_feat(87), I3 =>  inp_feat(509), I4 =>  inp_feat(290), I5 =>  inp_feat(74), I6 =>  inp_feat(250), I7 =>  inp_feat(235)); 
C_40_S_0_L_2_inst : LUT8 generic map(INIT => "0000100010001010100010001000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100011101000100010000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_0_L_2_out, I0 =>  inp_feat(183), I1 =>  inp_feat(407), I2 =>  inp_feat(475), I3 =>  inp_feat(415), I4 =>  inp_feat(73), I5 =>  inp_feat(81), I6 =>  inp_feat(116), I7 =>  inp_feat(211)); 
C_40_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000001000100000001100100000000000000000000000100011001000100010000101000010000000100011001000000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_0_L_3_out, I0 =>  inp_feat(4), I1 =>  inp_feat(38), I2 =>  inp_feat(351), I3 =>  inp_feat(73), I4 =>  inp_feat(20), I5 =>  inp_feat(504), I6 =>  inp_feat(316), I7 =>  inp_feat(251)); 
C_40_S_0_L_4_inst : LUT8 generic map(INIT => "0000000001110100010101010101010000000000000000000001010100000000000000000000000000010100000000010000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000") port map( O =>C_40_S_0_L_4_out, I0 =>  inp_feat(484), I1 =>  inp_feat(402), I2 =>  inp_feat(298), I3 =>  inp_feat(410), I4 =>  inp_feat(316), I5 =>  inp_feat(446), I6 =>  inp_feat(116), I7 =>  inp_feat(287)); 
C_40_S_0_L_5_inst : LUT8 generic map(INIT => "0010000011110000101000000000000000000000010100000010000011000000000000000000000000000000000000000000000000000000000000000000000010100011001000000000000000100000011110111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000") port map( O =>C_40_S_0_L_5_out, I0 =>  inp_feat(457), I1 =>  inp_feat(73), I2 =>  inp_feat(336), I3 =>  inp_feat(384), I4 =>  inp_feat(151), I5 =>  inp_feat(505), I6 =>  inp_feat(294), I7 =>  inp_feat(364)); 
C_40_S_0_L_6_inst : LUT8 generic map(INIT => "1011001110010001011100000001000100000001000100000000000000000000100000000000000000000000000000000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_0_L_6_out, I0 =>  inp_feat(471), I1 =>  inp_feat(452), I2 =>  inp_feat(133), I3 =>  inp_feat(264), I4 =>  inp_feat(486), I5 =>  inp_feat(116), I6 =>  inp_feat(287), I7 =>  inp_feat(251)); 
C_40_S_0_L_7_inst : LUT8 generic map(INIT => "0000000011000000000000000000000000010010001000000000000000000010000000000000000000000000000000000000000000000000000000000000000011110001111100000101000110000000101100101111000000010001100000000000000000010000000000000000000000000000000000010000000100000000") port map( O =>C_40_S_0_L_7_out, I0 =>  inp_feat(376), I1 =>  inp_feat(384), I2 =>  inp_feat(201), I3 =>  inp_feat(75), I4 =>  inp_feat(302), I5 =>  inp_feat(249), I6 =>  inp_feat(296), I7 =>  inp_feat(452)); 
C_40_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000011011000000000000000000000011000000100000000000000000000000001010100000000000000000000000001000100010000000000000000000000000000000000000000000000000000010110000001000000000000000000000000000000000000000000000000000001010001000100000000000000000") port map( O =>C_40_S_1_L_0_out, I0 =>  inp_feat(229), I1 =>  inp_feat(73), I2 =>  inp_feat(448), I3 =>  inp_feat(315), I4 =>  inp_feat(499), I5 =>  inp_feat(109), I6 =>  inp_feat(2), I7 =>  inp_feat(74)); 
C_40_S_1_L_1_inst : LUT8 generic map(INIT => "0011111111111100000001010000111000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_1_L_1_out, I0 =>  inp_feat(73), I1 =>  inp_feat(115), I2 =>  inp_feat(40), I3 =>  inp_feat(351), I4 =>  inp_feat(504), I5 =>  inp_feat(251), I6 =>  inp_feat(68), I7 =>  inp_feat(416)); 
C_40_S_1_L_2_inst : LUT8 generic map(INIT => "1000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000011100000100000001100100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_1_L_2_out, I0 =>  inp_feat(354), I1 =>  inp_feat(407), I2 =>  inp_feat(287), I3 =>  inp_feat(469), I4 =>  inp_feat(388), I5 =>  inp_feat(485), I6 =>  inp_feat(87), I7 =>  inp_feat(204)); 
C_40_S_1_L_3_inst : LUT8 generic map(INIT => "1001010011000100000100001000000000000000100000000000000010000000000000000000000000100000000000000000000000000000000000001000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_1_L_3_out, I0 =>  inp_feat(166), I1 =>  inp_feat(252), I2 =>  inp_feat(84), I3 =>  inp_feat(431), I4 =>  inp_feat(360), I5 =>  inp_feat(408), I6 =>  inp_feat(296), I7 =>  inp_feat(29)); 
C_40_S_1_L_4_inst : LUT8 generic map(INIT => "1000110000000100000000000000000000001000101010000000000000000000100011101000100000001000000000001000000010001000000000000000000000000000000000000000000000000000000000001010000000000000000000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_1_L_4_out, I0 =>  inp_feat(29), I1 =>  inp_feat(407), I2 =>  inp_feat(384), I3 =>  inp_feat(1), I4 =>  inp_feat(183), I5 =>  inp_feat(31), I6 =>  inp_feat(452), I7 =>  inp_feat(362)); 
C_40_S_1_L_5_inst : LUT8 generic map(INIT => "0101000000000000011001000000000000000000000000000011000000000000010010010000000000000010000000000000000000000000000000000000000011110000000000000011000000000000000000000000000000100000000000000111010000010000000000000000000001001000000000000000000000000000") port map( O =>C_40_S_1_L_5_out, I0 =>  inp_feat(328), I1 =>  inp_feat(448), I2 =>  inp_feat(398), I3 =>  inp_feat(336), I4 =>  inp_feat(31), I5 =>  inp_feat(446), I6 =>  inp_feat(285), I7 =>  inp_feat(273)); 
C_40_S_1_L_6_inst : LUT8 generic map(INIT => "1101010000000000010101011101000000010000000001000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_1_L_6_out, I0 =>  inp_feat(484), I1 =>  inp_feat(50), I2 =>  inp_feat(296), I3 =>  inp_feat(486), I4 =>  inp_feat(17), I5 =>  inp_feat(446), I6 =>  inp_feat(259), I7 =>  inp_feat(87)); 
C_40_S_1_L_7_inst : LUT8 generic map(INIT => "1001100000010000000000000000000001000001000000000000000000000000101000100000000010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_1_L_7_out, I0 =>  inp_feat(151), I1 =>  inp_feat(77), I2 =>  inp_feat(504), I3 =>  inp_feat(290), I4 =>  inp_feat(81), I5 =>  inp_feat(485), I6 =>  inp_feat(380), I7 =>  inp_feat(469)); 
C_40_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_0_out, I0 =>  inp_feat(287), I1 =>  inp_feat(5), I2 =>  inp_feat(290), I3 =>  inp_feat(130), I4 =>  inp_feat(179), I5 =>  inp_feat(241), I6 =>  inp_feat(251), I7 =>  inp_feat(92)); 
C_40_S_2_L_1_inst : LUT8 generic map(INIT => "0001000011110100000000000000000001110010001100000000000000000000011101001111000000000000000000001101000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_1_out, I0 =>  inp_feat(328), I1 =>  inp_feat(1), I2 =>  inp_feat(354), I3 =>  inp_feat(402), I4 =>  inp_feat(87), I5 =>  inp_feat(480), I6 =>  inp_feat(52), I7 =>  inp_feat(362)); 
C_40_S_2_L_2_inst : LUT8 generic map(INIT => "0001011100000000000011110000010110001100000011001101110100010000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_2_out, I0 =>  inp_feat(283), I1 =>  inp_feat(504), I2 =>  inp_feat(419), I3 =>  inp_feat(407), I4 =>  inp_feat(480), I5 =>  inp_feat(52), I6 =>  inp_feat(362), I7 =>  inp_feat(357)); 
C_40_S_2_L_3_inst : LUT8 generic map(INIT => "0000000010101000110001001100100000000000100000001000100010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_3_out, I0 =>  inp_feat(359), I1 =>  inp_feat(34), I2 =>  inp_feat(387), I3 =>  inp_feat(410), I4 =>  inp_feat(316), I5 =>  inp_feat(179), I6 =>  inp_feat(446), I7 =>  inp_feat(132)); 
C_40_S_2_L_4_inst : LUT8 generic map(INIT => "1110001000000000001000100000000011101110000010001000000000000000000000000000000000000000000000001000100000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_4_out, I0 =>  inp_feat(336), I1 =>  inp_feat(248), I2 =>  inp_feat(115), I3 =>  inp_feat(29), I4 =>  inp_feat(446), I5 =>  inp_feat(134), I6 =>  inp_feat(97), I7 =>  inp_feat(251)); 
C_40_S_2_L_5_inst : LUT8 generic map(INIT => "0010000001100111000000000111101101100010000001000010100000101100000000000000001100000000000000010011000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_5_out, I0 =>  inp_feat(445), I1 =>  inp_feat(73), I2 =>  inp_feat(248), I3 =>  inp_feat(1), I4 =>  inp_feat(31), I5 =>  inp_feat(504), I6 =>  inp_feat(127), I7 =>  inp_feat(469)); 
C_40_S_2_L_6_inst : LUT8 generic map(INIT => "0110101010001010001010110000101001011010110011010000001000000000000000000000000000000000100000000000000000001001000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_6_out, I0 =>  inp_feat(398), I1 =>  inp_feat(161), I2 =>  inp_feat(273), I3 =>  inp_feat(20), I4 =>  inp_feat(318), I5 =>  inp_feat(285), I6 =>  inp_feat(407), I7 =>  inp_feat(469)); 
C_40_S_2_L_7_inst : LUT8 generic map(INIT => "0001000011000000100100000010000011000000000000001111000000000000000000000000000000000000010000000100010001010000010100010001010110000000000000000000000000100100000000010001000000000000000000000000000100000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_2_L_7_out, I0 =>  inp_feat(92), I1 =>  inp_feat(274), I2 =>  inp_feat(183), I3 =>  inp_feat(93), I4 =>  inp_feat(420), I5 =>  inp_feat(50), I6 =>  inp_feat(341), I7 =>  inp_feat(296)); 
C_40_S_3_L_0_inst : LUT8 generic map(INIT => "0001000100000000010000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000100100000011100000010000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_40_S_3_L_0_out, I0 =>  inp_feat(134), I1 =>  inp_feat(339), I2 =>  inp_feat(367), I3 =>  inp_feat(302), I4 =>  inp_feat(247), I5 =>  inp_feat(51), I6 =>  inp_feat(251), I7 =>  inp_feat(92)); 
C_40_S_3_L_1_inst : LUT8 generic map(INIT => "1000000011110110000000001010000011100000110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_3_L_1_out, I0 =>  inp_feat(201), I1 =>  inp_feat(126), I2 =>  inp_feat(116), I3 =>  inp_feat(20), I4 =>  inp_feat(362), I5 =>  inp_feat(425), I6 =>  inp_feat(87), I7 =>  inp_feat(68)); 
C_40_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000101000000000000010001000000000000000000000000000000000000000001000000000000000000000000000000010111010100000000001001000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_3_L_2_out, I0 =>  inp_feat(354), I1 =>  inp_feat(226), I2 =>  inp_feat(493), I3 =>  inp_feat(29), I4 =>  inp_feat(407), I5 =>  inp_feat(152), I6 =>  inp_feat(287), I7 =>  inp_feat(452)); 
C_40_S_3_L_3_inst : LUT8 generic map(INIT => "0000010100001010000000001010001000000001000010000000000010000000001010100000100000101010000000101000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_40_S_3_L_3_out, I0 =>  inp_feat(308), I1 =>  inp_feat(20), I2 =>  inp_feat(1), I3 =>  inp_feat(384), I4 =>  inp_feat(505), I5 =>  inp_feat(504), I6 =>  inp_feat(73), I7 =>  inp_feat(100)); 
C_40_S_3_L_4_inst : LUT8 generic map(INIT => "1000001010100010101000001010101100000000100010001000000000001000000000100010000000000011100000001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_3_L_4_out, I0 =>  inp_feat(4), I1 =>  inp_feat(351), I2 =>  inp_feat(364), I3 =>  inp_feat(478), I4 =>  inp_feat(71), I5 =>  inp_feat(509), I6 =>  inp_feat(458), I7 =>  inp_feat(100)); 
C_40_S_3_L_5_inst : LUT8 generic map(INIT => "0001000001110000000000000000000000000000000100000000000010000000110100000101000001000000100000001000000001010100100000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000") port map( O =>C_40_S_3_L_5_out, I0 =>  inp_feat(221), I1 =>  inp_feat(31), I2 =>  inp_feat(29), I3 =>  inp_feat(249), I4 =>  inp_feat(309), I5 =>  inp_feat(17), I6 =>  inp_feat(273), I7 =>  inp_feat(362)); 
C_40_S_3_L_6_inst : LUT8 generic map(INIT => "1100110000000000010011100000001001111101000000100010101000001000010000100000000000001000000000000000000000000000001000100000001000000100000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_3_L_6_out, I0 =>  inp_feat(221), I1 =>  inp_feat(242), I2 =>  inp_feat(273), I3 =>  inp_feat(290), I4 =>  inp_feat(490), I5 =>  inp_feat(157), I6 =>  inp_feat(296), I7 =>  inp_feat(171)); 
C_40_S_3_L_7_inst : LUT8 generic map(INIT => "0001110100000000101001000010000000010011000000000000100000000000000001000000000010011100000000001111101000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_40_S_3_L_7_out, I0 =>  inp_feat(99), I1 =>  inp_feat(115), I2 =>  inp_feat(402), I3 =>  inp_feat(172), I4 =>  inp_feat(248), I5 =>  inp_feat(195), I6 =>  inp_feat(50), I7 =>  inp_feat(251)); 
C_40_S_4_L_0_inst : LUT8 generic map(INIT => "0000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010100010000000000000011000000010000000101000000000000000000000000000000000000000000000000000001000000000000000000000000000000") port map( O =>C_40_S_4_L_0_out, I0 =>  inp_feat(484), I1 =>  inp_feat(260), I2 =>  inp_feat(487), I3 =>  inp_feat(402), I4 =>  inp_feat(23), I5 =>  inp_feat(395), I6 =>  inp_feat(353), I7 =>  inp_feat(316)); 
C_40_S_4_L_1_inst : LUT8 generic map(INIT => "1100011100000100111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000110001000100100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_4_L_1_out, I0 =>  inp_feat(204), I1 =>  inp_feat(71), I2 =>  inp_feat(402), I3 =>  inp_feat(162), I4 =>  inp_feat(505), I5 =>  inp_feat(289), I6 =>  inp_feat(362), I7 =>  inp_feat(157)); 
C_40_S_4_L_2_inst : LUT8 generic map(INIT => "1000000000001010000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000101000000000000010101000101010100000000000001000100010101011101000000000000000000010000010000000000000000000000010000000001000000000000000000000") port map( O =>C_40_S_4_L_2_out, I0 =>  inp_feat(87), I1 =>  inp_feat(494), I2 =>  inp_feat(46), I3 =>  inp_feat(134), I4 =>  inp_feat(119), I5 =>  inp_feat(301), I6 =>  inp_feat(446), I7 =>  inp_feat(452)); 
C_40_S_4_L_3_inst : LUT8 generic map(INIT => "0000000010010001000000000000000000000000101001000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000010000000000000000000000001011110100000000000001000000000000000000000000000000000000000000000100110000000000000000") port map( O =>C_40_S_4_L_3_out, I0 =>  inp_feat(154), I1 =>  inp_feat(201), I2 =>  inp_feat(274), I3 =>  inp_feat(452), I4 =>  inp_feat(287), I5 =>  inp_feat(331), I6 =>  inp_feat(290), I7 =>  inp_feat(298)); 
C_40_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000011000000010001000000000001000000111000001100010000000000000001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_4_L_4_out, I0 =>  inp_feat(171), I1 =>  inp_feat(296), I2 =>  inp_feat(403), I3 =>  inp_feat(504), I4 =>  inp_feat(469), I5 =>  inp_feat(452), I6 =>  inp_feat(182), I7 =>  inp_feat(221)); 
C_40_S_4_L_5_inst : LUT8 generic map(INIT => "0010101100000000000000101000000000000000000000000000100000000000101010100000100000110000000010000101100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000001000000000000000000000000000") port map( O =>C_40_S_4_L_5_out, I0 =>  inp_feat(387), I1 =>  inp_feat(445), I2 =>  inp_feat(115), I3 =>  inp_feat(335), I4 =>  inp_feat(302), I5 =>  inp_feat(29), I6 =>  inp_feat(20), I7 =>  inp_feat(289)); 
C_40_S_4_L_6_inst : LUT8 generic map(INIT => "1001001010010000000000000000100010111010100010000000000010000000001100010110000100000000000000001111111110010000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000") port map( O =>C_40_S_4_L_6_out, I0 =>  inp_feat(262), I1 =>  inp_feat(384), I2 =>  inp_feat(71), I3 =>  inp_feat(285), I4 =>  inp_feat(100), I5 =>  inp_feat(73), I6 =>  inp_feat(249), I7 =>  inp_feat(163)); 
C_40_S_4_L_7_inst : LUT8 generic map(INIT => "0000000011000000000000000000000010001010001000001010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010000010100000001000000010100010100000000000000000000000000000") port map( O =>C_40_S_4_L_7_out, I0 =>  inp_feat(287), I1 =>  inp_feat(464), I2 =>  inp_feat(407), I3 =>  inp_feat(171), I4 =>  inp_feat(444), I5 =>  inp_feat(134), I6 =>  inp_feat(1), I7 =>  inp_feat(109)); 
C_41_S_0_L_0_inst : LUT8 generic map(INIT => "1111101111111111110110001111101111101110001000001100100010000000001011100000100110001010101010110000000000000000100010001000000010101000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_41_S_0_L_0_out, I0 =>  inp_feat(266), I1 =>  inp_feat(232), I2 =>  inp_feat(183), I3 =>  inp_feat(3), I4 =>  inp_feat(34), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_41_S_0_L_1_inst : LUT8 generic map(INIT => "0111111100010100111111110100111100001100000000000010000001000000101101011000011110110111110001011010010111000001000000110000000110110000000001001010000000000000100010000000000000000000000000001000100000000100100000000000000000000000000000000000000000000000") port map( O =>C_41_S_0_L_1_out, I0 =>  inp_feat(80), I1 =>  inp_feat(209), I2 =>  inp_feat(281), I3 =>  inp_feat(109), I4 =>  inp_feat(437), I5 =>  inp_feat(448), I6 =>  inp_feat(287), I7 =>  inp_feat(132)); 
C_41_S_0_L_2_inst : LUT8 generic map(INIT => "1100010010100000101011001110100011001100111000101110111011100100110010001000000011001000110010000100000010000000110010001100000000000000001000101000000011000100100001001111001011101100111011001100000000000000110000000000000000000000000000000000000000000000") port map( O =>C_41_S_0_L_2_out, I0 =>  inp_feat(471), I1 =>  inp_feat(301), I2 =>  inp_feat(410), I3 =>  inp_feat(339), I4 =>  inp_feat(387), I5 =>  inp_feat(222), I6 =>  inp_feat(123), I7 =>  inp_feat(452)); 
C_41_S_0_L_3_inst : LUT8 generic map(INIT => "1100110001001100111111011011010110101100000011000000000000000000111011000000110000000000000000001100110000001100000000000000000000001100000000001000000000000000010011000000000000000000000000001010100000000000100000000000000010000100000000000000000000000000") port map( O =>C_41_S_0_L_3_out, I0 =>  inp_feat(151), I1 =>  inp_feat(73), I2 =>  inp_feat(34), I3 =>  inp_feat(402), I4 =>  inp_feat(28), I5 =>  inp_feat(509), I6 =>  inp_feat(495), I7 =>  inp_feat(419)); 
C_41_S_0_L_4_inst : LUT8 generic map(INIT => "1111110001000101011110000100000101101100000001000000000000000000111100001000000011010000100001000110000000000000000000000000000011001101110001001111110010001101110011000000010001000000000000001100000000000000110100000000100001000000000000001100000000000000") port map( O =>C_41_S_0_L_4_out, I0 =>  inp_feat(444), I1 =>  inp_feat(464), I2 =>  inp_feat(381), I3 =>  inp_feat(134), I4 =>  inp_feat(239), I5 =>  inp_feat(1), I6 =>  inp_feat(29), I7 =>  inp_feat(290)); 
C_41_S_0_L_5_inst : LUT8 generic map(INIT => "0101010111010000011100010101000010111010011000001010001010000000101000001000000010000000000000000010001100100000111000000010000010110011000000000011001000100000101110001010001000110010001000001000000000000000001000000000000010110000101000000011000000100000") port map( O =>C_41_S_0_L_5_out, I0 =>  inp_feat(409), I1 =>  inp_feat(154), I2 =>  inp_feat(179), I3 =>  inp_feat(480), I4 =>  inp_feat(109), I5 =>  inp_feat(19), I6 =>  inp_feat(504), I7 =>  inp_feat(29)); 
C_41_S_0_L_6_inst : LUT8 generic map(INIT => "0101110111000000100011100000001011111101000000001010101000000000011111110100000001000000000000001101110101000000011010100100000000001101110011001100010001001101100011000000000010000000000000000101010100000000100000000000000000000000010000000111000000000000") port map( O =>C_41_S_0_L_6_out, I0 =>  inp_feat(336), I1 =>  inp_feat(504), I2 =>  inp_feat(407), I3 =>  inp_feat(137), I4 =>  inp_feat(229), I5 =>  inp_feat(388), I6 =>  inp_feat(390), I7 =>  inp_feat(41)); 
C_41_S_0_L_7_inst : LUT8 generic map(INIT => "0001001011011001110000110100000011011101110100010000000000000000110010111101010111001111110010011101110101010101010000000000000010100000000000000000000000000000101010000000000000000000000000001000100000000000100000000000000000001000000010000000000000000000") port map( O =>C_41_S_0_L_7_out, I0 =>  inp_feat(448), I1 =>  inp_feat(242), I2 =>  inp_feat(221), I3 =>  inp_feat(207), I4 =>  inp_feat(470), I5 =>  inp_feat(87), I6 =>  inp_feat(172), I7 =>  inp_feat(438)); 
C_41_S_1_L_0_inst : LUT8 generic map(INIT => "0101110011011100110011001000000011101110111011100010000000000000111011001111111011001100111000001010111010101110100000001010001000000010011010100000000010100000000010100000000000000000000000000000011001100010010000001010001000000010001000100000001000100000") port map( O =>C_41_S_1_L_0_out, I0 =>  inp_feat(222), I1 =>  inp_feat(284), I2 =>  inp_feat(409), I3 =>  inp_feat(229), I4 =>  inp_feat(364), I5 =>  inp_feat(401), I6 =>  inp_feat(437), I7 =>  inp_feat(179)); 
C_41_S_1_L_1_inst : LUT8 generic map(INIT => "0101110111010101101000000000000011010000110100000101000011100000011000000000000011100000001000000111000011010000111100001001000010100000111000001010000011000000000000001100000001000000111000001111000011110000110010010110000001000000110000001101000011000000") port map( O =>C_41_S_1_L_1_out, I0 =>  inp_feat(87), I1 =>  inp_feat(88), I2 =>  inp_feat(199), I3 =>  inp_feat(221), I4 =>  inp_feat(37), I5 =>  inp_feat(387), I6 =>  inp_feat(52), I7 =>  inp_feat(81)); 
C_41_S_1_L_2_inst : LUT8 generic map(INIT => "1111101010000000111100101000000010111010000000001011000000000000111100001000000011111000100000001010101100000000111111111000000010111000101000100011000000000000100000101111101001000000110000011000000010100000101100000000000011000000110100001111000111010011") port map( O =>C_41_S_1_L_2_out, I0 =>  inp_feat(329), I1 =>  inp_feat(302), I2 =>  inp_feat(134), I3 =>  inp_feat(493), I4 =>  inp_feat(130), I5 =>  inp_feat(467), I6 =>  inp_feat(81), I7 =>  inp_feat(274)); 
C_41_S_1_L_3_inst : LUT8 generic map(INIT => "1100100011100001101000101011110111110000001000001000000010000000100000000000000010000000000000001111000000000000000000000000000010100000000000001010000010000000100100001000000010001000100010000000000000000000000000000000100000000000100000000000000010000000") port map( O =>C_41_S_1_L_3_out, I0 =>  inp_feat(73), I1 =>  inp_feat(376), I2 =>  inp_feat(179), I3 =>  inp_feat(19), I4 =>  inp_feat(29), I5 =>  inp_feat(160), I6 =>  inp_feat(1), I7 =>  inp_feat(446)); 
C_41_S_1_L_4_inst : LUT8 generic map(INIT => "1010001010000000111000011100000010010000100000001000000000000000111111110000000011010101110000011111111100000000110111011000001011110000100000001111000010000000100000001000000010100000100000001111110000000000000000000000000000000000000000000000000000000000") port map( O =>C_41_S_1_L_4_out, I0 =>  inp_feat(41), I1 =>  inp_feat(509), I2 =>  inp_feat(20), I3 =>  inp_feat(1), I4 =>  inp_feat(178), I5 =>  inp_feat(109), I6 =>  inp_feat(446), I7 =>  inp_feat(232)); 
C_41_S_1_L_5_inst : LUT8 generic map(INIT => "1101100001010000011000000000000011110111000000001011000000000000100100000000000011111000000000000001110000000000110110000000000011101111110010001100011100000000111011110000000011111111000000001100000010000000100010000000000011001100000000001000100000000000") port map( O =>C_41_S_1_L_5_out, I0 =>  inp_feat(290), I1 =>  inp_feat(445), I2 =>  inp_feat(402), I3 =>  inp_feat(152), I4 =>  inp_feat(211), I5 =>  inp_feat(296), I6 =>  inp_feat(229), I7 =>  inp_feat(388)); 
C_41_S_1_L_6_inst : LUT8 generic map(INIT => "1110110110001000100011000000100010001111000010000000000000000000110011000100000001001100000000001100010110001000000001000000000011101100000010000000000000000000100001110000101000001000000000001100111000000000100011000000000011001101000011011100101000001000") port map( O =>C_41_S_1_L_6_out, I0 =>  inp_feat(460), I1 =>  inp_feat(199), I2 =>  inp_feat(336), I3 =>  inp_feat(134), I4 =>  inp_feat(73), I5 =>  inp_feat(478), I6 =>  inp_feat(340), I7 =>  inp_feat(461)); 
C_41_S_1_L_7_inst : LUT8 generic map(INIT => "1110101001001000010010001100010001001010111100000000000011110000110011001111110011000100111110001100000011110000000000001111000011101100111000001010000011100000101000001010000010100000101000001100000011000000010000001100010010000000000000000000000000000000") port map( O =>C_41_S_1_L_7_out, I0 =>  inp_feat(493), I1 =>  inp_feat(378), I2 =>  inp_feat(167), I3 =>  inp_feat(232), I4 =>  inp_feat(439), I5 =>  inp_feat(132), I6 =>  inp_feat(494), I7 =>  inp_feat(401)); 
C_41_S_2_L_0_inst : LUT8 generic map(INIT => "1010101011001000101011111111111110101010100000001010000000001000110111001111110010111011111111111000000010001000000000001010101000101010100000000010100000001010101010101000000010101010100000000010100010001000000000001000001000101000101010000000100010100000") port map( O =>C_41_S_2_L_0_out, I0 =>  inp_feat(235), I1 =>  inp_feat(340), I2 =>  inp_feat(383), I3 =>  inp_feat(388), I4 =>  inp_feat(41), I5 =>  inp_feat(80), I6 =>  inp_feat(296), I7 =>  inp_feat(109)); 
C_41_S_2_L_1_inst : LUT8 generic map(INIT => "1011011100100000110101011101010110000011000000000001000000010101101110110111001111110000111101011000000000000000010100000101000110110010100000101100000000000000000000000000000000000000000000000110000000100000110000001010000000000000000000000010000000000000") port map( O =>C_41_S_2_L_1_out, I0 =>  inp_feat(40), I1 =>  inp_feat(407), I2 =>  inp_feat(273), I3 =>  inp_feat(92), I4 =>  inp_feat(438), I5 =>  inp_feat(133), I6 =>  inp_feat(5), I7 =>  inp_feat(380)); 
C_41_S_2_L_2_inst : LUT8 generic map(INIT => "0100100011101100100000000010000010001100101010001000100010000000110100100010111101100011111110101111111011111010101010001010001011100000100010000000000000000000111100001010000000000000000000001010000010000000000000000000000011000000000000000000000000000000") port map( O =>C_41_S_2_L_2_out, I0 =>  inp_feat(504), I1 =>  inp_feat(509), I2 =>  inp_feat(109), I3 =>  inp_feat(362), I4 =>  inp_feat(92), I5 =>  inp_feat(232), I6 =>  inp_feat(437), I7 =>  inp_feat(132)); 
C_41_S_2_L_3_inst : LUT8 generic map(INIT => "1111010101000011111100001111001011101100110001000010000000000000111000001110000011110000010000001110000001000000101000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000011000000000000000100000000000000010000000000000") port map( O =>C_41_S_2_L_3_out, I0 =>  inp_feat(387), I1 =>  inp_feat(7), I2 =>  inp_feat(410), I3 =>  inp_feat(402), I4 =>  inp_feat(431), I5 =>  inp_feat(495), I6 =>  inp_feat(437), I7 =>  inp_feat(202)); 
C_41_S_2_L_4_inst : LUT8 generic map(INIT => "0000100000101010000111110000000011100010101010101101011100000000000000000000101000000001000000001000000010101010100000010000000010001010000010101000101000000010110000000000000010000000000000000000000000000000000000000000000011000000000000000000000000000000") port map( O =>C_41_S_2_L_4_out, I0 =>  inp_feat(278), I1 =>  inp_feat(431), I2 =>  inp_feat(232), I3 =>  inp_feat(28), I4 =>  inp_feat(509), I5 =>  inp_feat(357), I6 =>  inp_feat(73), I7 =>  inp_feat(495)); 
C_41_S_2_L_5_inst : LUT8 generic map(INIT => "0001111001100010100011110000011011100111000101101010111000001111111110000001000011001111000010000100110100000000000011110000101010110110001111111100001001001011001000010011011011101111010011111110111001111110010010110000111101100111000001010010011100001110") port map( O =>C_41_S_2_L_5_out, I0 =>  inp_feat(41), I1 =>  inp_feat(121), I2 =>  inp_feat(167), I3 =>  inp_feat(461), I4 =>  inp_feat(80), I5 =>  inp_feat(281), I6 =>  inp_feat(88), I7 =>  inp_feat(307)); 
C_41_S_2_L_6_inst : LUT8 generic map(INIT => "0000110111110000100100011011000001010001110101000000000000100000111111111000000011110001101000000000000000000000100000000010000010010100110110000111000011110011011010011111111001000000110100001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_41_S_2_L_6_out, I0 =>  inp_feat(290), I1 =>  inp_feat(448), I2 =>  inp_feat(504), I3 =>  inp_feat(172), I4 =>  inp_feat(256), I5 =>  inp_feat(115), I6 =>  inp_feat(253), I7 =>  inp_feat(336)); 
C_41_S_2_L_7_inst : LUT8 generic map(INIT => "1110111010001011101110000011001010001000100010101101000000000000100011000000000000110000111100000000000000000000000000000000000001000000000000001011000000000000100000000000000011110000000000000000000000100000001000000000000000000000000000000000000000000000") port map( O =>C_41_S_2_L_7_out, I0 =>  inp_feat(115), I1 =>  inp_feat(178), I2 =>  inp_feat(68), I3 =>  inp_feat(121), I4 =>  inp_feat(19), I5 =>  inp_feat(504), I6 =>  inp_feat(137), I7 =>  inp_feat(92)); 
C_41_S_3_L_0_inst : LUT8 generic map(INIT => "0111111110101000100010101010101100001010000000000000100010000000001011101010000010001000001010100000001000000000000010000000000010101100100010001000100010100000010011000000100010001000100000000000100010000000100010001010100000001000000000001000000010000000") port map( O =>C_41_S_3_L_0_out, I0 =>  inp_feat(134), I1 =>  inp_feat(29), I2 =>  inp_feat(336), I3 =>  inp_feat(450), I4 =>  inp_feat(232), I5 =>  inp_feat(109), I6 =>  inp_feat(88), I7 =>  inp_feat(281)); 
C_41_S_3_L_1_inst : LUT8 generic map(INIT => "0100100111100011111010001110100000100000000000101100101011000000110010000000101110001000100010100000000000000000001010101000101000000100010101000100000000100000000000000000000000000000000000000101010011011101100010001000000000000000000000000000000000000000") port map( O =>C_41_S_3_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(448), I2 =>  inp_feat(93), I3 =>  inp_feat(387), I4 =>  inp_feat(302), I5 =>  inp_feat(432), I6 =>  inp_feat(253), I7 =>  inp_feat(452)); 
C_41_S_3_L_2_inst : LUT8 generic map(INIT => "0111110111111000001100010100000010110011110111000001000000000000101000001110100001000000010000001000000010000000000000000000000000010000101010000101000001010000110000001100110000000000000000000000000001000000000000000000000001000000010000000000000000000000") port map( O =>C_41_S_3_L_2_out, I0 =>  inp_feat(154), I1 =>  inp_feat(81), I2 =>  inp_feat(410), I3 =>  inp_feat(388), I4 =>  inp_feat(115), I5 =>  inp_feat(253), I6 =>  inp_feat(192), I7 =>  inp_feat(92)); 
C_41_S_3_L_3_inst : LUT8 generic map(INIT => "1100001010000010110001001010111011011011111110111111111010001000100011101010111111001100110011101010110010111111010011001101101011011000000000011011010111010000111010111011101100011000101000011010111010001101110111011100110110101111101111110000110111111111") port map( O =>C_41_S_3_L_3_out, I0 =>  inp_feat(383), I1 =>  inp_feat(109), I2 =>  inp_feat(307), I3 =>  inp_feat(409), I4 =>  inp_feat(41), I5 =>  inp_feat(80), I6 =>  inp_feat(388), I7 =>  inp_feat(238)); 
C_41_S_3_L_4_inst : LUT8 generic map(INIT => "1001001011101010101000001110000010101010100000000000000010000010101100001000000001110010101100101000000010000000000000001010000011111000101010100000000010100010101010001010000000000010101000100000000000000010000000000010000010000010101000101000000010100010") port map( O =>C_41_S_3_L_4_out, I0 =>  inp_feat(73), I1 =>  inp_feat(7), I2 =>  inp_feat(204), I3 =>  inp_feat(302), I4 =>  inp_feat(15), I5 =>  inp_feat(253), I6 =>  inp_feat(242), I7 =>  inp_feat(388)); 
C_41_S_3_L_5_inst : LUT8 generic map(INIT => "0111001110000100110100001101010011110001110000000111000001010000001010100010000000000000100000000100001000000000000000001100000010101011101010101100000110100000101100000010000000000000101100000000000000000000000000000000000000100000000000000000000000000000") port map( O =>C_41_S_3_L_5_out, I0 =>  inp_feat(162), I1 =>  inp_feat(428), I2 =>  inp_feat(134), I3 =>  inp_feat(29), I4 =>  inp_feat(228), I5 =>  inp_feat(88), I6 =>  inp_feat(419), I7 =>  inp_feat(207)); 
C_41_S_3_L_6_inst : LUT8 generic map(INIT => "0011101111000100000000001000000011001100110000001001111010001000100010000100110000100000000010001100110011001100101010100100100010000000001010000000000010001010100010001000100000000000000010001000000010000000000000000000100000000000100010000000000000000000") port map( O =>C_41_S_3_L_6_out, I0 =>  inp_feat(504), I1 =>  inp_feat(36), I2 =>  inp_feat(431), I3 =>  inp_feat(80), I4 =>  inp_feat(461), I5 =>  inp_feat(372), I6 =>  inp_feat(229), I7 =>  inp_feat(76)); 
C_41_S_3_L_7_inst : LUT8 generic map(INIT => "0010011110010010010101010100000000000011111010100001100110001011100101111011101100100000000000100011001100111011001010110011001111111111010001001010011100000000000110101000100000001010101010101100010000001110000000000000000000000000000010000000000010000000") port map( O =>C_41_S_3_L_7_out, I0 =>  inp_feat(310), I1 =>  inp_feat(183), I2 =>  inp_feat(154), I3 =>  inp_feat(444), I4 =>  inp_feat(298), I5 =>  inp_feat(438), I6 =>  inp_feat(446), I7 =>  inp_feat(11)); 
C_41_S_4_L_0_inst : LUT8 generic map(INIT => "0101010111011100110000001111010111101110010101010100010001000100011111101111111001011000111101011111111000001110010101000101010011011000101111110000100010100101010111000101010101000000000001001000100011101110110001011110010111010101010111000101010001010101") port map( O =>C_41_S_4_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(109), I2 =>  inp_feat(121), I3 =>  inp_feat(80), I4 =>  inp_feat(461), I5 =>  inp_feat(88), I6 =>  inp_feat(307), I7 =>  inp_feat(238)); 
C_41_S_4_L_1_inst : LUT8 generic map(INIT => "0010001010101000111010101100010010101000101000101110111111000010110011111010000010101010000000001101111100100010001000100000000010000000000010001100110011000000000010100000000011000100110001000000100000000000000000000000000010000010000000000000000000000000") port map( O =>C_41_S_4_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(448), I2 =>  inp_feat(290), I3 =>  inp_feat(130), I4 =>  inp_feat(444), I5 =>  inp_feat(11), I6 =>  inp_feat(296), I7 =>  inp_feat(255)); 
C_41_S_4_L_2_inst : LUT8 generic map(INIT => "1011101011111010101110001011001011111010111100101110001010101010111010001100000000000000000000001100110010000000110001000000000010100001101001100000001000101000100000101000100011001010000000101010100000001110000000000000101011001000000000001100110000000000") port map( O =>C_41_S_4_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(307), I2 =>  inp_feat(364), I3 =>  inp_feat(232), I4 =>  inp_feat(88), I5 =>  inp_feat(437), I6 =>  inp_feat(182), I7 =>  inp_feat(340)); 
C_41_S_4_L_3_inst : LUT8 generic map(INIT => "0011110111101111101111101000111100100000000000000000000000000000101111110001101010101111110111110010000010000000000000001000100010000000000000001000000000000000110000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_41_S_4_L_3_out, I0 =>  inp_feat(36), I1 =>  inp_feat(207), I2 =>  inp_feat(217), I3 =>  inp_feat(140), I4 =>  inp_feat(444), I5 =>  inp_feat(288), I6 =>  inp_feat(73), I7 =>  inp_feat(495)); 
C_41_S_4_L_4_inst : LUT8 generic map(INIT => "0000110001001010111010100000111001111000100000001111000000000000000000001000000010000000000000001000100010000000100000000000000010101010101011101000100011111110101000001000000010100000000000001000000010000000000000000000000010000000100000000000000000000000") port map( O =>C_41_S_4_L_4_out, I0 =>  inp_feat(152), I1 =>  inp_feat(497), I2 =>  inp_feat(140), I3 =>  inp_feat(60), I4 =>  inp_feat(130), I5 =>  inp_feat(388), I6 =>  inp_feat(253), I7 =>  inp_feat(408)); 
C_41_S_4_L_5_inst : LUT8 generic map(INIT => "1111101010100000111011110000000001101010000000100000000000000000100100111011100011111011000010100111000100010000100000000000000011100100010000001111000010110000100000000000000011110000001000000100000000110000101100001000000000000000000000000000000000000000") port map( O =>C_41_S_4_L_5_out, I0 =>  inp_feat(373), I1 =>  inp_feat(302), I2 =>  inp_feat(228), I3 =>  inp_feat(134), I4 =>  inp_feat(68), I5 =>  inp_feat(484), I6 =>  inp_feat(41), I7 =>  inp_feat(281)); 
C_41_S_4_L_6_inst : LUT8 generic map(INIT => "1110010111110101111010101111001000000000110000001000101011010010111111011111011100100000001000100101000100000000000100010000000011000000110000001010000011110000010000001100000000000000111100000000000000000000100000000000000000000000000000000001000100000000") port map( O =>C_41_S_4_L_6_out, I0 =>  inp_feat(287), I1 =>  inp_feat(387), I2 =>  inp_feat(402), I3 =>  inp_feat(339), I4 =>  inp_feat(289), I5 =>  inp_feat(1), I6 =>  inp_feat(296), I7 =>  inp_feat(109)); 
C_41_S_4_L_7_inst : LUT8 generic map(INIT => "0111001111010111000010000100000011010111110001111000100000000000000010100000000000001000100000001010001000000000000010001000000010111010110000000000000010000000100000001000000010001000100010000000000000000000100000001000000000000000000000001000100010001000") port map( O =>C_41_S_4_L_7_out, I0 =>  inp_feat(446), I1 =>  inp_feat(287), I2 =>  inp_feat(372), I3 =>  inp_feat(383), I4 =>  inp_feat(489), I5 =>  inp_feat(388), I6 =>  inp_feat(431), I7 =>  inp_feat(495)); 
C_42_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000001000100010110000100000000010000000100000000000000000000010100000101010000000000010001000000000000000000000000010000000000000000000100000001000001010000000000000000000000000000000000000000000001000100000000000100010") port map( O =>C_42_S_0_L_0_out, I0 =>  inp_feat(29), I1 =>  inp_feat(202), I2 =>  inp_feat(204), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_42_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000100000011100000010000001010000000000000000000000000000000000000000000000000000001000000000000000000000011000000010100000100111001010000010000001100000010000000000000000100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_0_L_1_out, I0 =>  inp_feat(452), I1 =>  inp_feat(407), I2 =>  inp_feat(336), I3 =>  inp_feat(384), I4 =>  inp_feat(509), I5 =>  inp_feat(1), I6 =>  inp_feat(408), I7 =>  inp_feat(273)); 
C_42_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000110010000010001000000000000000000000000000000000000000101100001010001010000000101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_0_L_2_out, I0 =>  inp_feat(81), I1 =>  inp_feat(504), I2 =>  inp_feat(130), I3 =>  inp_feat(378), I4 =>  inp_feat(320), I5 =>  inp_feat(487), I6 =>  inp_feat(204), I7 =>  inp_feat(251)); 
C_42_S_0_L_3_inst : LUT8 generic map(INIT => "0001000000000000000000000010000000000000000000000000000000000000000000000000000001100000000000000010000000000000000000000011001011110000000000001111000100000000000100000001000000010000000000000000000000000000001000000000000000000000000000000010000000000010") port map( O =>C_42_S_0_L_3_out, I0 =>  inp_feat(316), I1 =>  inp_feat(40), I2 =>  inp_feat(274), I3 =>  inp_feat(6), I4 =>  inp_feat(285), I5 =>  inp_feat(497), I6 =>  inp_feat(19), I7 =>  inp_feat(179)); 
C_42_S_0_L_4_inst : LUT8 generic map(INIT => "0001000011110000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000100010000000000000000000100000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_0_L_4_out, I0 =>  inp_feat(497), I1 =>  inp_feat(411), I2 =>  inp_feat(159), I3 =>  inp_feat(178), I4 =>  inp_feat(487), I5 =>  inp_feat(154), I6 =>  inp_feat(183), I7 =>  inp_feat(20)); 
C_42_S_0_L_5_inst : LUT8 generic map(INIT => "1000000010100000000000000000000011000000100010000000100000000000000000001000000000000000000000001100110011101100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000") port map( O =>C_42_S_0_L_5_out, I0 =>  inp_feat(407), I1 =>  inp_feat(469), I2 =>  inp_feat(455), I3 =>  inp_feat(473), I4 =>  inp_feat(183), I5 =>  inp_feat(204), I6 =>  inp_feat(222), I7 =>  inp_feat(84)); 
C_42_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000101000001000000000000000000000000000000000001000100000000010000010000000011000100000000000000000000000000000001010101010001000000010000000000000000000000000000000000000000000001000000000000000001010101010101000000000000000000000000000101000") port map( O =>C_42_S_0_L_6_out, I0 =>  inp_feat(19), I1 =>  inp_feat(302), I2 =>  inp_feat(347), I3 =>  inp_feat(420), I4 =>  inp_feat(273), I5 =>  inp_feat(388), I6 =>  inp_feat(285), I7 =>  inp_feat(286)); 
C_42_S_0_L_7_inst : LUT8 generic map(INIT => "1110000011010000010000000100100000000000111100000000000010001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_0_L_7_out, I0 =>  inp_feat(445), I1 =>  inp_feat(411), I2 =>  inp_feat(84), I3 =>  inp_feat(221), I4 =>  inp_feat(20), I5 =>  inp_feat(504), I6 =>  inp_feat(241), I7 =>  inp_feat(158)); 
C_42_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000001000100010110000100000000010000000100000000000000000000010100000101010000000000010001000000000000000000000000010000000000000000000100000001000001010000000000000000000000000000000000000000000001000100000000000100010") port map( O =>C_42_S_1_L_0_out, I0 =>  inp_feat(29), I1 =>  inp_feat(202), I2 =>  inp_feat(204), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_42_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000100000000000000010100000000000001000000000000000000000000000000000000000000000000000000000000000001000001010000000010001000000001010100110000000100000000000000010100000000000000000000000000000000000010001000000000000000000000000000000000000") port map( O =>C_42_S_1_L_1_out, I0 =>  inp_feat(413), I1 =>  inp_feat(504), I2 =>  inp_feat(403), I3 =>  inp_feat(296), I4 =>  inp_feat(452), I5 =>  inp_feat(1), I6 =>  inp_feat(408), I7 =>  inp_feat(273)); 
C_42_S_1_L_2_inst : LUT8 generic map(INIT => "0000001000010110000001000000111000000000000000000000000000000010111111001110110001001100001011100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_1_L_2_out, I0 =>  inp_feat(402), I1 =>  inp_feat(77), I2 =>  inp_feat(288), I3 =>  inp_feat(378), I4 =>  inp_feat(317), I5 =>  inp_feat(469), I6 =>  inp_feat(445), I7 =>  inp_feat(487)); 
C_42_S_1_L_3_inst : LUT8 generic map(INIT => "0000000011000000000001000100000110100000101000000000000000000000111000001000000000000000011110000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_1_L_3_out, I0 =>  inp_feat(352), I1 =>  inp_feat(139), I2 =>  inp_feat(469), I3 =>  inp_feat(445), I4 =>  inp_feat(158), I5 =>  inp_feat(2), I6 =>  inp_feat(204), I7 =>  inp_feat(183)); 
C_42_S_1_L_4_inst : LUT8 generic map(INIT => "0000001100000000000100000000000010110011000000100000000000000000101010000000100100000000000000001010101000001010000010000000000000000000000000000000000000000000100010000000000000000000000000000001100000000000000000000000000010001000000000000000000000000000") port map( O =>C_42_S_1_L_4_out, I0 =>  inp_feat(373), I1 =>  inp_feat(472), I2 =>  inp_feat(420), I3 =>  inp_feat(407), I4 =>  inp_feat(183), I5 =>  inp_feat(445), I6 =>  inp_feat(92), I7 =>  inp_feat(154)); 
C_42_S_1_L_5_inst : LUT8 generic map(INIT => "1000000000001000000000000000000001001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001010000000000000100110000001100110000000000100010000000000000000000000000000000000000000000000000000000000000010001") port map( O =>C_42_S_1_L_5_out, I0 =>  inp_feat(41), I1 =>  inp_feat(84), I2 =>  inp_feat(504), I3 =>  inp_feat(283), I4 =>  inp_feat(81), I5 =>  inp_feat(109), I6 =>  inp_feat(383), I7 =>  inp_feat(247)); 
C_42_S_1_L_6_inst : LUT8 generic map(INIT => "1100000000000000000000000000000010000100100010000000000000000000111000001111000101100000001000001010010010100000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_1_L_6_out, I0 =>  inp_feat(151), I1 =>  inp_feat(154), I2 =>  inp_feat(29), I3 =>  inp_feat(458), I4 =>  inp_feat(274), I5 =>  inp_feat(301), I6 =>  inp_feat(20), I7 =>  inp_feat(487)); 
C_42_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000100010000000000000000000000000000000000000000000000000000000000010111000000000100000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000100011101010000000000000000000000000000000100000000010100000") port map( O =>C_42_S_1_L_7_out, I0 =>  inp_feat(469), I1 =>  inp_feat(179), I2 =>  inp_feat(199), I3 =>  inp_feat(221), I4 =>  inp_feat(488), I5 =>  inp_feat(119), I6 =>  inp_feat(247), I7 =>  inp_feat(364)); 
C_42_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000001000100010110000100000000010000000100000000000000000000010100000101010000000000010001000000000000000000000000010000000000000000000100000001000001010000000000000000000000000000000000000000000001000100000000000100010") port map( O =>C_42_S_2_L_0_out, I0 =>  inp_feat(29), I1 =>  inp_feat(202), I2 =>  inp_feat(204), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_42_S_2_L_1_inst : LUT8 generic map(INIT => "1100010100000100000000000000000000000000000000000000000000000000110111010000010000100010000000000100000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000") port map( O =>C_42_S_2_L_1_out, I0 =>  inp_feat(484), I1 =>  inp_feat(229), I2 =>  inp_feat(199), I3 =>  inp_feat(251), I4 =>  inp_feat(413), I5 =>  inp_feat(116), I6 =>  inp_feat(273), I7 =>  inp_feat(408)); 
C_42_S_2_L_2_inst : LUT8 generic map(INIT => "0000001000000000000000000000000000010111001000110000000100000000111101010000010000000000000000001111111100000101000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_2_L_2_out, I0 =>  inp_feat(52), I1 =>  inp_feat(152), I2 =>  inp_feat(301), I3 =>  inp_feat(407), I4 =>  inp_feat(469), I5 =>  inp_feat(247), I6 =>  inp_feat(452), I7 =>  inp_feat(487)); 
C_42_S_2_L_3_inst : LUT8 generic map(INIT => "0000010000001100000000000000000000000000000011000000000000000000010011001100110000000000000000000000110011001100000000000000000000000000000000000000000000000000010000000001000000000000000000000000010011000000000000000000000000000000110000000000000000000000") port map( O =>C_42_S_2_L_3_out, I0 =>  inp_feat(211), I1 =>  inp_feat(485), I2 =>  inp_feat(73), I3 =>  inp_feat(415), I4 =>  inp_feat(183), I5 =>  inp_feat(445), I6 =>  inp_feat(204), I7 =>  inp_feat(284)); 
C_42_S_2_L_4_inst : LUT8 generic map(INIT => "1101100000010001010000000001000000000000000000010000000100000000110011001100110100000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_2_L_4_out, I0 =>  inp_feat(450), I1 =>  inp_feat(27), I2 =>  inp_feat(412), I3 =>  inp_feat(411), I4 =>  inp_feat(436), I5 =>  inp_feat(469), I6 =>  inp_feat(179), I7 =>  inp_feat(154)); 
C_42_S_2_L_5_inst : LUT8 generic map(INIT => "1011001010110001000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000011000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_2_L_5_out, I0 =>  inp_feat(222), I1 =>  inp_feat(298), I2 =>  inp_feat(129), I3 =>  inp_feat(244), I4 =>  inp_feat(256), I5 =>  inp_feat(217), I6 =>  inp_feat(487), I7 =>  inp_feat(428)); 
C_42_S_2_L_6_inst : LUT8 generic map(INIT => "0000001000000000001000110000000000000000000000000000000000000010001000100000000000100010000000000000000000000000000000000000000000000010000000000000101000000000000000000000000000000000000000000010101100000000000000100000000000000000000000000000000000000000") port map( O =>C_42_S_2_L_6_out, I0 =>  inp_feat(183), I1 =>  inp_feat(316), I2 =>  inp_feat(58), I3 =>  inp_feat(172), I4 =>  inp_feat(31), I5 =>  inp_feat(407), I6 =>  inp_feat(273), I7 =>  inp_feat(402)); 
C_42_S_2_L_7_inst : LUT8 generic map(INIT => "0000011010001000000000000000000000000000000000000000000010000000000011111100100100000000000000000000010000000000000000000000000000000100000000100000000010101000000000000000000000000000000000000000111100001000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_2_L_7_out, I0 =>  inp_feat(170), I1 =>  inp_feat(154), I2 =>  inp_feat(415), I3 =>  inp_feat(221), I4 =>  inp_feat(238), I5 =>  inp_feat(183), I6 =>  inp_feat(445), I7 =>  inp_feat(314)); 
C_42_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000001000100010110000100000000010000000100000000000000000000010100000101010000000000010001000000000000000000000000010000000000000000000100000001000001010000000000000000000000000000000000000000000001000100000000000100010") port map( O =>C_42_S_3_L_0_out, I0 =>  inp_feat(29), I1 =>  inp_feat(202), I2 =>  inp_feat(204), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_42_S_3_L_1_inst : LUT8 generic map(INIT => "1011100010111011000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_3_L_1_out, I0 =>  inp_feat(357), I1 =>  inp_feat(221), I2 =>  inp_feat(274), I3 =>  inp_feat(445), I4 =>  inp_feat(124), I5 =>  inp_feat(251), I6 =>  inp_feat(338), I7 =>  inp_feat(408)); 
C_42_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000010000000100000001000000001000000110010001000000000000000000000000000100000000000000000000000000000000000000000000000000000001100001010001000011011010000010010001000101010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_3_L_2_out, I0 =>  inp_feat(242), I1 =>  inp_feat(222), I2 =>  inp_feat(445), I3 =>  inp_feat(58), I4 =>  inp_feat(221), I5 =>  inp_feat(415), I6 =>  inp_feat(487), I7 =>  inp_feat(273)); 
C_42_S_3_L_3_inst : LUT8 generic map(INIT => "0000001010001000000000100000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100010100000000000000000000000001000000000000000000000001010000010100010000000000000000000000000100010000000100000001000") port map( O =>C_42_S_3_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(291), I2 =>  inp_feat(301), I3 =>  inp_feat(415), I4 =>  inp_feat(302), I5 =>  inp_feat(193), I6 =>  inp_feat(364), I7 =>  inp_feat(1)); 
C_42_S_3_L_4_inst : LUT8 generic map(INIT => "0111110000101100000000001000000001001100000000000100110001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_3_L_4_out, I0 =>  inp_feat(445), I1 =>  inp_feat(148), I2 =>  inp_feat(302), I3 =>  inp_feat(383), I4 =>  inp_feat(354), I5 =>  inp_feat(98), I6 =>  inp_feat(487), I7 =>  inp_feat(469)); 
C_42_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000100000001000000000000000110011110000000000000000000000001010010010100000101010100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000110000000000000") port map( O =>C_42_S_3_L_5_out, I0 =>  inp_feat(157), I1 =>  inp_feat(264), I2 =>  inp_feat(274), I3 =>  inp_feat(81), I4 =>  inp_feat(6), I5 =>  inp_feat(247), I6 =>  inp_feat(273), I7 =>  inp_feat(407)); 
C_42_S_3_L_6_inst : LUT8 generic map(INIT => "0000000110010011110100001111000000000001000000000100000000000001000000000000000000000000100000000000000000000000000000000000000000000000001000001000000010110000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_42_S_3_L_6_out, I0 =>  inp_feat(504), I1 =>  inp_feat(229), I2 =>  inp_feat(336), I3 =>  inp_feat(412), I4 =>  inp_feat(316), I5 =>  inp_feat(407), I6 =>  inp_feat(388), I7 =>  inp_feat(112)); 
C_42_S_3_L_7_inst : LUT8 generic map(INIT => "0001000101011101000000001000000000000000000000000000100000000000001011010101110100001000100000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000") port map( O =>C_42_S_3_L_7_out, I0 =>  inp_feat(291), I1 =>  inp_feat(71), I2 =>  inp_feat(187), I3 =>  inp_feat(452), I4 =>  inp_feat(475), I5 =>  inp_feat(81), I6 =>  inp_feat(161), I7 =>  inp_feat(486)); 
C_42_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000001000100010110000100000000010000000100000000000000000000010100000101010000000000010001000000000000000000000000010000000000000000000100000001000001010000000000000000000000000000000000000000000001000100000000000100010") port map( O =>C_42_S_4_L_0_out, I0 =>  inp_feat(29), I1 =>  inp_feat(202), I2 =>  inp_feat(204), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_42_S_4_L_1_inst : LUT8 generic map(INIT => "1011100010111011000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_4_L_1_out, I0 =>  inp_feat(357), I1 =>  inp_feat(221), I2 =>  inp_feat(274), I3 =>  inp_feat(445), I4 =>  inp_feat(124), I5 =>  inp_feat(251), I6 =>  inp_feat(338), I7 =>  inp_feat(408)); 
C_42_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000010000000100000001000000001000000110010001000000000000000000000000000100000000000000000000000000000000000000000000000000000001100001010001000011011010000010010001000101010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_4_L_2_out, I0 =>  inp_feat(242), I1 =>  inp_feat(222), I2 =>  inp_feat(445), I3 =>  inp_feat(58), I4 =>  inp_feat(221), I5 =>  inp_feat(415), I6 =>  inp_feat(487), I7 =>  inp_feat(273)); 
C_42_S_4_L_3_inst : LUT8 generic map(INIT => "0000001010001000000000100000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100010100000000000000000000000001000000000000000000000001010000010100010000000000000000000000000100010000000100000001000") port map( O =>C_42_S_4_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(291), I2 =>  inp_feat(301), I3 =>  inp_feat(415), I4 =>  inp_feat(302), I5 =>  inp_feat(193), I6 =>  inp_feat(364), I7 =>  inp_feat(1)); 
C_42_S_4_L_4_inst : LUT8 generic map(INIT => "0111110000101100000000001000000001001100000000000100110001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_4_L_4_out, I0 =>  inp_feat(445), I1 =>  inp_feat(148), I2 =>  inp_feat(302), I3 =>  inp_feat(383), I4 =>  inp_feat(354), I5 =>  inp_feat(98), I6 =>  inp_feat(487), I7 =>  inp_feat(469)); 
C_42_S_4_L_5_inst : LUT8 generic map(INIT => "0000001100000000000000000000000000000110011011110000000000000000101100110000011000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000010001000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_4_L_5_out, I0 =>  inp_feat(384), I1 =>  inp_feat(204), I2 =>  inp_feat(179), I3 =>  inp_feat(109), I4 =>  inp_feat(289), I5 =>  inp_feat(1), I6 =>  inp_feat(376), I7 =>  inp_feat(407)); 
C_42_S_4_L_6_inst : LUT8 generic map(INIT => "0000000010000000110000000000101001000000100000001101100010001100000000000000000000000000000000000000100000000000011000000000000000000000000000000000000000000000000000001000000011000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_4_L_6_out, I0 =>  inp_feat(274), I1 =>  inp_feat(387), I2 =>  inp_feat(229), I3 =>  inp_feat(247), I4 =>  inp_feat(273), I5 =>  inp_feat(484), I6 =>  inp_feat(183), I7 =>  inp_feat(438)); 
C_42_S_4_L_7_inst : LUT8 generic map(INIT => "0010001000100000001000000000000000000000000000000000000000000000001000001010000000000000000000001000000010000000000000001000000010000000101000100010000010100000000000000000000010000000101000000000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_42_S_4_L_7_out, I0 =>  inp_feat(383), I1 =>  inp_feat(328), I2 =>  inp_feat(274), I3 =>  inp_feat(218), I4 =>  inp_feat(117), I5 =>  inp_feat(256), I6 =>  inp_feat(439), I7 =>  inp_feat(412)); 
C_43_S_0_L_0_inst : LUT8 generic map(INIT => "1111111111111111100010001000100011111001111100001111100111000000101000101000000000000000000000000000000110100000000000000000000010001000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_43_S_0_L_0_out, I0 =>  inp_feat(329), I1 =>  inp_feat(469), I2 =>  inp_feat(78), I3 =>  inp_feat(362), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_43_S_0_L_1_inst : LUT8 generic map(INIT => "1100111011101111100011101110111010001010101010101000001000000010111011001010001010000000001000101000000010101010101010001010101000001000000000000000000000000000001000000000000000000000000000001100010000000000000000000000000000000000000000000000000000000000") port map( O =>C_43_S_0_L_1_out, I0 =>  inp_feat(134), I1 =>  inp_feat(31), I2 =>  inp_feat(290), I3 =>  inp_feat(413), I4 =>  inp_feat(448), I5 =>  inp_feat(504), I6 =>  inp_feat(250), I7 =>  inp_feat(235)); 
C_43_S_0_L_2_inst : LUT8 generic map(INIT => "1110101111101010111110101010101110000000000010001110001010101010111011111010000010100000001000001000000000000000000000000000000000101000010000001010000011110100000000000000000010000000010000001011101010100000101000001010000000000000000000000000000000000000") port map( O =>C_43_S_0_L_2_out, I0 =>  inp_feat(179), I1 =>  inp_feat(166), I2 =>  inp_feat(288), I3 =>  inp_feat(411), I4 =>  inp_feat(29), I5 =>  inp_feat(425), I6 =>  inp_feat(87), I7 =>  inp_feat(273)); 
C_43_S_0_L_3_inst : LUT8 generic map(INIT => "0111111010101010101000100000000010000010101010001010001000000000001100001000100000100010001010001000000010101000001010100010100000000100101000000010001000000000000000000000000000100010000000000000000010100000001010101010100000000000100000000010101010001000") port map( O =>C_43_S_0_L_3_out, I0 =>  inp_feat(284), I1 =>  inp_feat(172), I2 =>  inp_feat(359), I3 =>  inp_feat(407), I4 =>  inp_feat(354), I5 =>  inp_feat(287), I6 =>  inp_feat(90), I7 =>  inp_feat(251)); 
C_43_S_0_L_4_inst : LUT8 generic map(INIT => "1000100100000000000010000000000011101010000000001110100010000000101010100000000010100000000000001100000011000000110000000000000010110010111100001000101110100000111011100000000011001111100000000000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_43_S_0_L_4_out, I0 =>  inp_feat(504), I1 =>  inp_feat(457), I2 =>  inp_feat(274), I3 =>  inp_feat(1), I4 =>  inp_feat(301), I5 =>  inp_feat(81), I6 =>  inp_feat(446), I7 =>  inp_feat(129)); 
C_43_S_0_L_5_inst : LUT8 generic map(INIT => "1110111011000011111010100000011100100110000101010000000000000000000000000000111010001100100000000100000000000001000011000000000010101010001010101000000000000000000000100000001000000000000000000010011000001010110001000000000000001110000000101000110000000000") port map( O =>C_43_S_0_L_5_out, I0 =>  inp_feat(446), I1 =>  inp_feat(180), I2 =>  inp_feat(302), I3 =>  inp_feat(485), I4 =>  inp_feat(287), I5 =>  inp_feat(383), I6 =>  inp_feat(456), I7 =>  inp_feat(253)); 
C_43_S_0_L_6_inst : LUT8 generic map(INIT => "0010111000010001110011001010000100000000000000001100110010100110101011110011111110101010001010110000000000000000000000001010101011100000000000001100100000000000010000000000000001000000000000001111001000000000000000000000000000000000000000000000000000000000") port map( O =>C_43_S_0_L_6_out, I0 =>  inp_feat(134), I1 =>  inp_feat(130), I2 =>  inp_feat(6), I3 =>  inp_feat(247), I4 =>  inp_feat(407), I5 =>  inp_feat(140), I6 =>  inp_feat(81), I7 =>  inp_feat(12)); 
C_43_S_0_L_7_inst : LUT8 generic map(INIT => "0011000011110000100000001011000011101101110111001100110000000000110001001010100011101100101000001000100000001000000010000000100010110000101100000100000010100000000000001000000000000000000000001010000010101000101000001010000000001000000010000000000000000000") port map( O =>C_43_S_0_L_7_out, I0 =>  inp_feat(75), I1 =>  inp_feat(207), I2 =>  inp_feat(415), I3 =>  inp_feat(457), I4 =>  inp_feat(301), I5 =>  inp_feat(388), I6 =>  inp_feat(251), I7 =>  inp_feat(445)); 
C_43_S_1_L_0_inst : LUT8 generic map(INIT => "1111111000001010111110100000000011001110110000101010101000000000100011100000101110001010000010000000000000000000000010000000000000101000000000100110100000000000010000000000000010110000011100111011000000110011011010111011111100000000000100010111001100110011") port map( O =>C_43_S_1_L_0_out, I0 =>  inp_feat(273), I1 =>  inp_feat(388), I2 =>  inp_feat(272), I3 =>  inp_feat(92), I4 =>  inp_feat(287), I5 =>  inp_feat(87), I6 =>  inp_feat(446), I7 =>  inp_feat(320)); 
C_43_S_1_L_1_inst : LUT8 generic map(INIT => "0101010001011110111100001101110000100011111111111100100011001000000100001011000000000000111100001010000000000000000000000000000011110000100000001010100010001000100000001000000000000000000000001001000000000000000000000000000010100000000000000000000000000000") port map( O =>C_43_S_1_L_1_out, I0 =>  inp_feat(336), I1 =>  inp_feat(41), I2 =>  inp_feat(273), I3 =>  inp_feat(407), I4 =>  inp_feat(354), I5 =>  inp_feat(387), I6 =>  inp_feat(299), I7 =>  inp_feat(93)); 
C_43_S_1_L_2_inst : LUT8 generic map(INIT => "0010111011100000101010001000100011000100000001000100010001000000111101000100010011000000000000001100010000000000110000000100000011100100000000001000110010100000110000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000") port map( O =>C_43_S_1_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(452), I2 =>  inp_feat(406), I3 =>  inp_feat(134), I4 =>  inp_feat(72), I5 =>  inp_feat(299), I6 =>  inp_feat(93), I7 =>  inp_feat(251)); 
C_43_S_1_L_3_inst : LUT8 generic map(INIT => "1110000001100010111010001010001010000000000000001000100000001000111100001010001000000000101000101110100010100010100010001010100010101010101010101000111110101111001000000000000010001000000000001010000010100000100000000000000000100000101000001000100010001000") port map( O =>C_43_S_1_L_3_out, I0 =>  inp_feat(73), I1 =>  inp_feat(285), I2 =>  inp_feat(109), I3 =>  inp_feat(1), I4 =>  inp_feat(289), I5 =>  inp_feat(204), I6 =>  inp_feat(407), I7 =>  inp_feat(438)); 
C_43_S_1_L_4_inst : LUT8 generic map(INIT => "0000000011000111111100001111010100000010000000100000000011110010001000001100000000000001000100000000000000000000000000000001001111110111110011100101010101110111010001110000011101010111110111110010001000100000000000000010000100000000000000000000000000000001") port map( O =>C_43_S_1_L_4_out, I0 =>  inp_feat(287), I1 =>  inp_feat(154), I2 =>  inp_feat(204), I3 =>  inp_feat(444), I4 =>  inp_feat(438), I5 =>  inp_feat(353), I6 =>  inp_feat(133), I7 =>  inp_feat(201)); 
C_43_S_1_L_5_inst : LUT8 generic map(INIT => "0011101111111111100000111111110010001010111111000000000011111100101101100010001000000000000000000010101110011010000000000000000010111101111111011111110111111111111111011111110100111101111111010001100000000000000000010000000000001001000010000000000000011011") port map( O =>C_43_S_1_L_5_out, I0 =>  inp_feat(318), I1 =>  inp_feat(336), I2 =>  inp_feat(229), I3 =>  inp_feat(100), I4 =>  inp_feat(61), I5 =>  inp_feat(291), I6 =>  inp_feat(504), I7 =>  inp_feat(469)); 
C_43_S_1_L_6_inst : LUT8 generic map(INIT => "1111101011001101110110001101100000001000000001000000000001000000100000000100110100000000000000001100000010000101000000000000000011001100010010110100111011101010000000000000001000000000000000000000000001000100000000000000000000000000000000000000000000000000") port map( O =>C_43_S_1_L_6_out, I0 =>  inp_feat(435), I1 =>  inp_feat(92), I2 =>  inp_feat(438), I3 =>  inp_feat(86), I4 =>  inp_feat(391), I5 =>  inp_feat(133), I6 =>  inp_feat(17), I7 =>  inp_feat(424)); 
C_43_S_1_L_7_inst : LUT8 generic map(INIT => "0111111100101000000000100000001001110111000010100010001100000010101010100000000000000000000000001000010000000000000000000000000011111111001000001111010100100010101111110010101001011111000000101010101000100000101100010000000000000110001000000011000000000000") port map( O =>C_43_S_1_L_7_out, I0 =>  inp_feat(274), I1 =>  inp_feat(81), I2 =>  inp_feat(265), I3 =>  inp_feat(248), I4 =>  inp_feat(61), I5 =>  inp_feat(221), I6 =>  inp_feat(504), I7 =>  inp_feat(158)); 
C_43_S_2_L_0_inst : LUT8 generic map(INIT => "1111110011111110110000001100000010100000101110000000000000000000110000001111100000000000011000001111000011001100010010000000000000110000111011100000000011000000000000000000000000000000000000000000000011001010000000001100000000000000000000000000000000000000") port map( O =>C_43_S_2_L_0_out, I0 =>  inp_feat(431), I1 =>  inp_feat(204), I2 =>  inp_feat(262), I3 =>  inp_feat(86), I4 =>  inp_feat(73), I5 =>  inp_feat(356), I6 =>  inp_feat(61), I7 =>  inp_feat(251)); 
C_43_S_2_L_1_inst : LUT8 generic map(INIT => "0101110011110000100010000000000011001101000000001100110010000000110100010000000010000000000000000100000000000000010000000000000011001101100010001000000010000000010011010000000011001100000000001100110111001100100000001000000000000000000000000000000000000000") port map( O =>C_43_S_2_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(69), I2 =>  inp_feat(391), I3 =>  inp_feat(31), I4 =>  inp_feat(446), I5 =>  inp_feat(186), I6 =>  inp_feat(419), I7 =>  inp_feat(290)); 
C_43_S_2_L_2_inst : LUT8 generic map(INIT => "0000101010100011000001001100010010001010100000000000000011000000001111101100110110011111110011101000100010000000100000001100000011101110111111110000000000000000100010000000100000000000000000000000100000000000000000000000000000001000000000000000000000000000") port map( O =>C_43_S_2_L_2_out, I0 =>  inp_feat(471), I1 =>  inp_feat(410), I2 =>  inp_feat(25), I3 =>  inp_feat(201), I4 =>  inp_feat(94), I5 =>  inp_feat(100), I6 =>  inp_feat(108), I7 =>  inp_feat(423)); 
C_43_S_2_L_3_inst : LUT8 generic map(INIT => "1110010010101100111001001010110010101100111111010101110111111101111000000000100011001000011000001010100010001000111111101100110010101000100010001000000000000000000000000000100000000000000010000000000000001000000000000000000000000000000010000000100000001000") port map( O =>C_43_S_2_L_3_out, I0 =>  inp_feat(51), I1 =>  inp_feat(316), I2 =>  inp_feat(221), I3 =>  inp_feat(302), I4 =>  inp_feat(467), I5 =>  inp_feat(108), I6 =>  inp_feat(37), I7 =>  inp_feat(432)); 
C_43_S_2_L_4_inst : LUT8 generic map(INIT => "0111110101011111110001010000010111011111110101111100111100000101101100100000000000010000000000001000000000000000101000000000000011111101111100001101110101000100110100000101000011000100000000000000000000000000000000000000000010100000000000000010000000000000") port map( O =>C_43_S_2_L_4_out, I0 =>  inp_feat(336), I1 =>  inp_feat(88), I2 =>  inp_feat(81), I3 =>  inp_feat(504), I4 =>  inp_feat(301), I5 =>  inp_feat(362), I6 =>  inp_feat(112), I7 =>  inp_feat(87)); 
C_43_S_2_L_5_inst : LUT8 generic map(INIT => "0010011100000000111100000111000011001010000000001111110011110000111111110000001100110100010000001011111110010011111101011011010111101111000001000000000000000000010011000000000001000100000001000010011101000101010101010001010100000101000001010000010101000101") port map( O =>C_43_S_2_L_5_out, I0 =>  inp_feat(307), I1 =>  inp_feat(387), I2 =>  inp_feat(287), I3 =>  inp_feat(445), I4 =>  inp_feat(274), I5 =>  inp_feat(407), I6 =>  inp_feat(201), I7 =>  inp_feat(423)); 
C_43_S_2_L_6_inst : LUT8 generic map(INIT => "1111110011010001001111110111011111111000010110001111000000000000000010000001100101010100111111011000100011001000000000001000000000001000010000000000000000000000101000000100000001100000000000001000100000000000000000000000000010000000000000001000000010000000") port map( O =>C_43_S_2_L_6_out, I0 =>  inp_feat(287), I1 =>  inp_feat(353), I2 =>  inp_feat(486), I3 =>  inp_feat(296), I4 =>  inp_feat(239), I5 =>  inp_feat(108), I6 =>  inp_feat(274), I7 =>  inp_feat(247)); 
C_43_S_2_L_7_inst : LUT8 generic map(INIT => "1011111011100100000001001111010010000000110000000000000011100100101001000000000011110100111101001010000011000000001000000100000011100100100000000110010001000100100000000000000000000000010100001100110000100000110011000101110011000000000000000000000000000000") port map( O =>C_43_S_2_L_7_out, I0 =>  inp_feat(460), I1 =>  inp_feat(285), I2 =>  inp_feat(415), I3 =>  inp_feat(107), I4 =>  inp_feat(254), I5 =>  inp_feat(73), I6 =>  inp_feat(265), I7 =>  inp_feat(228)); 
C_43_S_3_L_0_inst : LUT8 generic map(INIT => "1111111100110111101000011011000111111111111100111001101000000000111011110000010110110000001000000100111101000000000000000000000000111111001100110011001100000001100001110000000110000010000000000000111100000000101100001011000000001111000000000000000000000000") port map( O =>C_43_S_3_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(494), I2 =>  inp_feat(121), I3 =>  inp_feat(484), I4 =>  inp_feat(134), I5 =>  inp_feat(265), I6 =>  inp_feat(251), I7 =>  inp_feat(61)); 
C_43_S_3_L_1_inst : LUT8 generic map(INIT => "0100110100001100111110010001000001100000000000001000000000000000110111011101010011110001110100000000000000000000000000000000000011111101110000001000100011000000110000000000000010000000000000001101110100000000100000000000000001010000000000000000000000000000") port map( O =>C_43_S_3_L_1_out, I0 =>  inp_feat(407), I1 =>  inp_feat(334), I2 =>  inp_feat(251), I3 =>  inp_feat(504), I4 =>  inp_feat(265), I5 =>  inp_feat(425), I6 =>  inp_feat(87), I7 =>  inp_feat(499)); 
C_43_S_3_L_2_inst : LUT8 generic map(INIT => "1111110111110000001110110011100011111111101100100010101000100010010100000001000000001001000110010011001100000001001100110000001110000111000000000000111100000010111011111010000000001111000000110000000000000000000000000000000000000001000000010000010000000000") port map( O =>C_43_S_3_L_2_out, I0 =>  inp_feat(494), I1 =>  inp_feat(4), I2 =>  inp_feat(364), I3 =>  inp_feat(504), I4 =>  inp_feat(408), I5 =>  inp_feat(336), I6 =>  inp_feat(419), I7 =>  inp_feat(273)); 
C_43_S_3_L_3_inst : LUT8 generic map(INIT => "0100101100001000100010000010000011111111110000101010001000000010110011001100110010000000000000001100000010000000000000000000000011000010011000100000000000000010010000100010001000000000000000000100000000000000000000000000000001000000000000000000000000000000") port map( O =>C_43_S_3_L_3_out, I0 =>  inp_feat(351), I1 =>  inp_feat(213), I2 =>  inp_feat(120), I3 =>  inp_feat(92), I4 =>  inp_feat(112), I5 =>  inp_feat(87), I6 =>  inp_feat(186), I7 =>  inp_feat(423)); 
C_43_S_3_L_4_inst : LUT8 generic map(INIT => "0100000111101000100010001010111110000000100010000000000010001000110000001100000000000000010001001101000011010000110001001100100011000000000000000000000000000000000000000000000000000000000000001101000001000001110000001100010011010000010100001100000011010001") port map( O =>C_43_S_3_L_4_out, I0 =>  inp_feat(469), I1 =>  inp_feat(179), I2 =>  inp_feat(152), I3 =>  inp_feat(336), I4 =>  inp_feat(84), I5 =>  inp_feat(465), I6 =>  inp_feat(48), I7 =>  inp_feat(37)); 
C_43_S_3_L_5_inst : LUT8 generic map(INIT => "1110110010001100110011001010110010100000101011101010000010101110000000001000000010000000100000000000000010001000100000000000000000100000000000001110000001100100001100011111111011000000111011100000000000000000100000000000000010010000101111111000000010000000") port map( O =>C_43_S_3_L_5_out, I0 =>  inp_feat(273), I1 =>  inp_feat(116), I2 =>  inp_feat(57), I3 =>  inp_feat(287), I4 =>  inp_feat(290), I5 =>  inp_feat(438), I6 =>  inp_feat(501), I7 =>  inp_feat(92)); 
C_43_S_3_L_6_inst : LUT8 generic map(INIT => "1010111000001000101110110001101110101100101011000010000000000000111010111000001111111011101110110000000000100000000000001010000001001111000011010000001100000011000011000100110000000000000000000000000100000011010000110000001100000000100000000000000010000000") port map( O =>C_43_S_3_L_6_out, I0 =>  inp_feat(328), I1 =>  inp_feat(364), I2 =>  inp_feat(407), I3 =>  inp_feat(221), I4 =>  inp_feat(408), I5 =>  inp_feat(327), I6 =>  inp_feat(265), I7 =>  inp_feat(251)); 
C_43_S_3_L_7_inst : LUT8 generic map(INIT => "1010000011111010010100001010000000111011101110100111000010010000110111110000001011010000000000001111001110000011101100000100000011101001111011111010000011001001111111111111111000010000111000001111111110001110111100001100000010110011000100101010000000000010") port map( O =>C_43_S_3_L_7_out, I0 =>  inp_feat(445), I1 =>  inp_feat(473), I2 =>  inp_feat(402), I3 =>  inp_feat(97), I4 =>  inp_feat(157), I5 =>  inp_feat(322), I6 =>  inp_feat(290), I7 =>  inp_feat(444)); 
C_43_S_4_L_0_inst : LUT8 generic map(INIT => "0100000111011000110011001000000001001100110011000000110101001100011011101000100010000000100000001111000010000000000000001100000011000111100110000000010000001100010001001000100000000100000011001111111110001000000000000000000011110000000010000000000000000000") port map( O =>C_43_S_4_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(92), I2 =>  inp_feat(108), I3 =>  inp_feat(100), I4 =>  inp_feat(37), I5 =>  inp_feat(48), I6 =>  inp_feat(347), I7 =>  inp_feat(5)); 
C_43_S_4_L_1_inst : LUT8 generic map(INIT => "0110101010101101011000101000000010100011101001111110101111000000101000001110101110000100111000001000001110100111001001001010000000000010000000111010101000000000000010110000000111001110000000000000000000000010010001000000000000000011000001110000000000000000") port map( O =>C_43_S_4_L_1_out, I0 =>  inp_feat(204), I1 =>  inp_feat(457), I2 =>  inp_feat(98), I3 =>  inp_feat(438), I4 =>  inp_feat(108), I5 =>  inp_feat(87), I6 =>  inp_feat(154), I7 =>  inp_feat(273)); 
C_43_S_4_L_2_inst : LUT8 generic map(INIT => "0101111101011000010111011000100011010101110110110000000010000000111111111001100110001000100010000011001110111011000000001000100011000000100000001000110000000000111000111111001100000000000000000010000000000010100010000000000000110011001100110000000000000000") port map( O =>C_43_S_4_L_2_out, I0 =>  inp_feat(362), I1 =>  inp_feat(262), I2 =>  inp_feat(274), I3 =>  inp_feat(464), I4 =>  inp_feat(450), I5 =>  inp_feat(500), I6 =>  inp_feat(296), I7 =>  inp_feat(251)); 
C_43_S_4_L_3_inst : LUT8 generic map(INIT => "1110110011100010110000001110000001110111110010101111011101011000111010100010001011110010100000001001000110101010111100000000001010101000001000000000000000100000011011110010101000100011101000100111001000100000000000000000001011111111001010100000001000100010") port map( O =>C_43_S_4_L_3_out, I0 =>  inp_feat(336), I1 =>  inp_feat(222), I2 =>  inp_feat(5), I3 =>  inp_feat(151), I4 =>  inp_feat(322), I5 =>  inp_feat(444), I6 =>  inp_feat(52), I7 =>  inp_feat(446)); 
C_43_S_4_L_4_inst : LUT8 generic map(INIT => "0111010001010001001100000101000011000000100000000000000000000000111110000111101111101000110100101000100001000000010000000000000001110101001100011111000010110000000000000001000000000000000000001110110101000001100010000000000000000000010000000000000000000000") port map( O =>C_43_S_4_L_4_out, I0 =>  inp_feat(108), I1 =>  inp_feat(336), I2 =>  inp_feat(204), I3 =>  inp_feat(301), I4 =>  inp_feat(134), I5 =>  inp_feat(117), I6 =>  inp_feat(494), I7 =>  inp_feat(154)); 
C_43_S_4_L_5_inst : LUT8 generic map(INIT => "0111111000101100101000101001001011011010001000001010100000101010001110100000000011110000000000001010000000000000001000000000000011101010001000001000000000000000101000101010000010000000000010001010101000000000000000000000000000100010000000000000000000000000") port map( O =>C_43_S_4_L_5_out, I0 =>  inp_feat(204), I1 =>  inp_feat(297), I2 =>  inp_feat(241), I3 =>  inp_feat(419), I4 =>  inp_feat(436), I5 =>  inp_feat(265), I6 =>  inp_feat(471), I7 =>  inp_feat(85)); 
C_43_S_4_L_6_inst : LUT8 generic map(INIT => "1111110010101000110000001000000011111101101000000000000000000000000000001000000000100000101000000010000010100000000000000000000011101111100010001100110010100000000101011000000000100000100000001000000010000000000000001000000010000000100000000000000010000000") port map( O =>C_43_S_4_L_6_out, I0 =>  inp_feat(309), I1 =>  inp_feat(88), I2 =>  inp_feat(439), I3 =>  inp_feat(68), I4 =>  inp_feat(397), I5 =>  inp_feat(391), I6 =>  inp_feat(14), I7 =>  inp_feat(265)); 
C_43_S_4_L_7_inst : LUT8 generic map(INIT => "1010001011101000111000111000100010001010000010001000100010001000010100000000000011111000100010000000000000001000000000001000000000000000110100001000100010001000000000000000100000000000100010001100000011001000110000001000100000000000100010001000000010001000") port map( O =>C_43_S_4_L_7_out, I0 =>  inp_feat(109), I1 =>  inp_feat(31), I2 =>  inp_feat(402), I3 =>  inp_feat(446), I4 =>  inp_feat(296), I5 =>  inp_feat(410), I6 =>  inp_feat(298), I7 =>  inp_feat(251)); 
C_44_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000001000000100000000000100000000000001000000000000000000000000000001100101111000000001010101000000000000000000000000000110000000000000010000000100000101000100000000000000000000000000000000000000000101010000000000010101010") port map( O =>C_44_S_0_L_0_out, I0 =>  inp_feat(260), I1 =>  inp_feat(412), I2 =>  inp_feat(480), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_44_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000001011101000000000111001000000000000000000000000000100000000000000000000000000000001100110000000000000000000000000000000000000000") port map( O =>C_44_S_0_L_1_out, I0 =>  inp_feat(134), I1 =>  inp_feat(419), I2 =>  inp_feat(270), I3 =>  inp_feat(335), I4 =>  inp_feat(109), I5 =>  inp_feat(251), I6 =>  inp_feat(74), I7 =>  inp_feat(235)); 
C_44_S_0_L_2_inst : LUT8 generic map(INIT => "1000000000100000101000000000000000000000000000000000000000000000111000001110000010000000000000001100000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_0_L_2_out, I0 =>  inp_feat(438), I1 =>  inp_feat(180), I2 =>  inp_feat(81), I3 =>  inp_feat(446), I4 =>  inp_feat(253), I5 =>  inp_feat(487), I6 =>  inp_feat(452), I7 =>  inp_feat(388)); 
C_44_S_0_L_3_inst : LUT8 generic map(INIT => "0011011100010111010101010101001100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101000000000101010100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_0_L_3_out, I0 =>  inp_feat(484), I1 =>  inp_feat(204), I2 =>  inp_feat(57), I3 =>  inp_feat(170), I4 =>  inp_feat(384), I5 =>  inp_feat(287), I6 =>  inp_feat(241), I7 =>  inp_feat(74)); 
C_44_S_0_L_4_inst : LUT8 generic map(INIT => "0111000001110011000100000110000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010110100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_0_L_4_out, I0 =>  inp_feat(484), I1 =>  inp_feat(204), I2 =>  inp_feat(171), I3 =>  inp_feat(134), I4 =>  inp_feat(201), I5 =>  inp_feat(388), I6 =>  inp_feat(241), I7 =>  inp_feat(169)); 
C_44_S_0_L_5_inst : LUT8 generic map(INIT => "0000101000000000100000000000000010001000100010010000000000000000000000010000000000000000000000001000100000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_0_L_5_out, I0 =>  inp_feat(94), I1 =>  inp_feat(158), I2 =>  inp_feat(57), I3 =>  inp_feat(407), I4 =>  inp_feat(287), I5 =>  inp_feat(92), I6 =>  inp_feat(242), I7 =>  inp_feat(438)); 
C_44_S_0_L_6_inst : LUT8 generic map(INIT => "1000000000001100000000000000000010100010101000000010000000000010000000000000000000000000000000000010000010000010000000000000000000000000000000000000000000000000100010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_0_L_6_out, I0 =>  inp_feat(34), I1 =>  inp_feat(381), I2 =>  inp_feat(383), I3 =>  inp_feat(154), I4 =>  inp_feat(290), I5 =>  inp_feat(40), I6 =>  inp_feat(388), I7 =>  inp_feat(438)); 
C_44_S_0_L_7_inst : LUT8 generic map(INIT => "0100000000000000000000000000000000000000100000000000000000000000010010000000100000000000000000000000100001111000000000000000000010000000000000000000000000000000110000001100000000000000000000001010000011000000000000000000000011000000111000000000000000000000") port map( O =>C_44_S_0_L_7_out, I0 =>  inp_feat(256), I1 =>  inp_feat(302), I2 =>  inp_feat(370), I3 =>  inp_feat(115), I4 =>  inp_feat(241), I5 =>  inp_feat(179), I6 =>  inp_feat(52), I7 =>  inp_feat(415)); 
C_44_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000001000000100000000000100000000000001000000000000000000000000000001100101111000000001010101000000000000000000000000000110000000000000010000000100000101000100000000000000000000000000000000000000000101010000000000010101010") port map( O =>C_44_S_1_L_0_out, I0 =>  inp_feat(260), I1 =>  inp_feat(412), I2 =>  inp_feat(480), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_44_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000001000000010000000000000000000000000000000000000000000000010000000000000001000100000000000000000000000000000000010110000001000001010000000100000000000000010000000000000000000000000000000100000000000000010000000000000000000000000000000000000") port map( O =>C_44_S_1_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(221), I2 =>  inp_feat(81), I3 =>  inp_feat(109), I4 =>  inp_feat(204), I5 =>  inp_feat(251), I6 =>  inp_feat(74), I7 =>  inp_feat(235)); 
C_44_S_1_L_2_inst : LUT8 generic map(INIT => "0010000000000000111000001000000000000000000000000000000000000000111100110101000010110000101100000001000010010000000000000010000000000000000000000000010000000000000000000000000000000000000000000001000100000000000100000001011000000000000000000000000000000000") port map( O =>C_44_S_1_L_2_out, I0 =>  inp_feat(420), I1 =>  inp_feat(92), I2 =>  inp_feat(171), I3 =>  inp_feat(201), I4 =>  inp_feat(402), I5 =>  inp_feat(487), I6 =>  inp_feat(452), I7 =>  inp_feat(388)); 
C_44_S_1_L_3_inst : LUT8 generic map(INIT => "0011101100001100001010110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000100010100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_1_L_3_out, I0 =>  inp_feat(388), I1 =>  inp_feat(402), I2 =>  inp_feat(452), I3 =>  inp_feat(183), I4 =>  inp_feat(201), I5 =>  inp_feat(411), I6 =>  inp_feat(241), I7 =>  inp_feat(179)); 
C_44_S_1_L_4_inst : LUT8 generic map(INIT => "0010111000001011001000101000001000100010001000100010001000000010000000001000100000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000") port map( O =>C_44_S_1_L_4_out, I0 =>  inp_feat(487), I1 =>  inp_feat(204), I2 =>  inp_feat(484), I3 =>  inp_feat(151), I4 =>  inp_feat(37), I5 =>  inp_feat(301), I6 =>  inp_feat(25), I7 =>  inp_feat(388)); 
C_44_S_1_L_5_inst : LUT8 generic map(INIT => "0110011100110011000100101111001100000010000000000000000000010000010100010000000010110000000100001000000000000000000100000001000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000") port map( O =>C_44_S_1_L_5_out, I0 =>  inp_feat(262), I1 =>  inp_feat(316), I2 =>  inp_feat(31), I3 =>  inp_feat(50), I4 =>  inp_feat(445), I5 =>  inp_feat(383), I6 =>  inp_feat(93), I7 =>  inp_feat(438)); 
C_44_S_1_L_6_inst : LUT8 generic map(INIT => "1100101010000000000000000000000000000000000000000000000000000000000010000001101000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_1_L_6_out, I0 =>  inp_feat(446), I1 =>  inp_feat(458), I2 =>  inp_feat(484), I3 =>  inp_feat(88), I4 =>  inp_feat(87), I5 =>  inp_feat(155), I6 =>  inp_feat(30), I7 =>  inp_feat(241)); 
C_44_S_1_L_7_inst : LUT8 generic map(INIT => "0010000000000010001010001000000000001000000010001000100000000000000000000000000010000000000000000000000000001000100010000000000000000000000000001100000000000000000000001100000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_44_S_1_L_7_out, I0 =>  inp_feat(407), I1 =>  inp_feat(296), I2 =>  inp_feat(402), I3 =>  inp_feat(446), I4 =>  inp_feat(57), I5 =>  inp_feat(442), I6 =>  inp_feat(438), I7 =>  inp_feat(236)); 
C_44_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000001000000100000000000100000000000001000000000000000000000000000001100101111000000001010101000000000000000000000000000110000000000000010000000100000101000100000000000000000000000000000000000000000101010000000000010101010") port map( O =>C_44_S_2_L_0_out, I0 =>  inp_feat(260), I1 =>  inp_feat(412), I2 =>  inp_feat(480), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_44_S_2_L_1_inst : LUT8 generic map(INIT => "1011001010101110000000100000001010000000111010100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_2_L_1_out, I0 =>  inp_feat(407), I1 =>  inp_feat(152), I2 =>  inp_feat(57), I3 =>  inp_feat(452), I4 =>  inp_feat(336), I5 =>  inp_feat(133), I6 =>  inp_feat(116), I7 =>  inp_feat(232)); 
C_44_S_2_L_2_inst : LUT8 generic map(INIT => "0101000001000000000000000000000011110000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000001010000000001000001000000000000111001001100010000000000100100010000000000000100000000000000000000000000000000000000000000000000") port map( O =>C_44_S_2_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(494), I2 =>  inp_feat(355), I3 =>  inp_feat(152), I4 =>  inp_feat(27), I5 =>  inp_feat(448), I6 =>  inp_feat(287), I7 =>  inp_feat(273)); 
C_44_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000001000000101001000000000000000000100000000100000000000000010000001000000011110111000000001000010000000000000000000000000000000000000000001000100000000000000000001010000010000000100000000000000000000100110000000000000000000000") port map( O =>C_44_S_2_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(154), I2 =>  inp_feat(157), I3 =>  inp_feat(235), I4 =>  inp_feat(183), I5 =>  inp_feat(134), I6 =>  inp_feat(316), I7 =>  inp_feat(419)); 
C_44_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000011110011000000010000000000000000000000000000000000000000000000000000000100000000000000000000000011001011000000000000000000000000111110000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_2_L_4_out, I0 =>  inp_feat(450), I1 =>  inp_feat(342), I2 =>  inp_feat(256), I3 =>  inp_feat(87), I4 =>  inp_feat(241), I5 =>  inp_feat(316), I6 =>  inp_feat(289), I7 =>  inp_feat(134)); 
C_44_S_2_L_5_inst : LUT8 generic map(INIT => "0101000001000000000000000000100000000000000000000000000000000000010000001110000010001000100000100000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000001000000000000000000000000000000000001000") port map( O =>C_44_S_2_L_5_out, I0 =>  inp_feat(202), I1 =>  inp_feat(487), I2 =>  inp_feat(486), I3 =>  inp_feat(204), I4 =>  inp_feat(242), I5 =>  inp_feat(388), I6 =>  inp_feat(134), I7 =>  inp_feat(438)); 
C_44_S_2_L_6_inst : LUT8 generic map(INIT => "0100001000010100000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_2_L_6_out, I0 =>  inp_feat(301), I1 =>  inp_feat(93), I2 =>  inp_feat(305), I3 =>  inp_feat(388), I4 =>  inp_feat(81), I5 =>  inp_feat(29), I6 =>  inp_feat(241), I7 =>  inp_feat(364)); 
C_44_S_2_L_7_inst : LUT8 generic map(INIT => "1100110000100100000000000000000010001110001000100000000000000000100001000000100000000000000000000000000000000000000000000000000001000000000010000000000000001000110000000000000000000000000000000000110000000100000000000000000000001100000000000000000000000000") port map( O =>C_44_S_2_L_7_out, I0 =>  inp_feat(420), I1 =>  inp_feat(81), I2 =>  inp_feat(52), I3 =>  inp_feat(383), I4 =>  inp_feat(34), I5 =>  inp_feat(444), I6 =>  inp_feat(201), I7 =>  inp_feat(93)); 
C_44_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000001000000100000000000100000000000001000000000000000000000000000001100101111000000001010101000000000000000000000000000110000000000000010000000100000101000100000000000000000000000000000000000000000101010000000000010101010") port map( O =>C_44_S_3_L_0_out, I0 =>  inp_feat(260), I1 =>  inp_feat(412), I2 =>  inp_feat(480), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_44_S_3_L_1_inst : LUT8 generic map(INIT => "1100010011010110000000000000001110000100110001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_3_L_1_out, I0 =>  inp_feat(316), I1 =>  inp_feat(370), I2 =>  inp_feat(36), I3 =>  inp_feat(61), I4 =>  inp_feat(336), I5 =>  inp_feat(133), I6 =>  inp_feat(116), I7 =>  inp_feat(232)); 
C_44_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000010000010000010100000000000110000001010101010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000010100000101000101010001010100010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_3_L_2_out, I0 =>  inp_feat(289), I1 =>  inp_feat(142), I2 =>  inp_feat(301), I3 =>  inp_feat(419), I4 =>  inp_feat(415), I5 =>  inp_feat(484), I6 =>  inp_feat(287), I7 =>  inp_feat(273)); 
C_44_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000010000110111000000000000000000011110000001001000000000000000000011000001010000000000000000000000000000100000000000000000000000000000000000100000000000000000000001000000000000000000000000000000010000000000000000000000000000") port map( O =>C_44_S_3_L_3_out, I0 =>  inp_feat(484), I1 =>  inp_feat(121), I2 =>  inp_feat(119), I3 =>  inp_feat(1), I4 =>  inp_feat(241), I5 =>  inp_feat(419), I6 =>  inp_feat(15), I7 =>  inp_feat(302)); 
C_44_S_3_L_4_inst : LUT8 generic map(INIT => "0001110010111000000000000000000000100000111111000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_3_L_4_out, I0 =>  inp_feat(108), I1 =>  inp_feat(152), I2 =>  inp_feat(157), I3 =>  inp_feat(484), I4 =>  inp_feat(241), I5 =>  inp_feat(419), I6 =>  inp_feat(81), I7 =>  inp_feat(251)); 
C_44_S_3_L_5_inst : LUT8 generic map(INIT => "0101000000000000010000000000000000010000010000000000000000000000111000001100000001000000000000000100010000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000100010000000000000000000100000001000000000000000000000000000000") port map( O =>C_44_S_3_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(334), I2 =>  inp_feat(487), I3 =>  inp_feat(486), I4 =>  inp_feat(388), I5 =>  inp_feat(446), I6 =>  inp_feat(134), I7 =>  inp_feat(438)); 
C_44_S_3_L_6_inst : LUT8 generic map(INIT => "1010000000000000001000000000000010101000001000001000000000000000000000001000000000000000000000000000000010100000000000000000000010100000100001000000000010000000000000101000000000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_3_L_6_out, I0 =>  inp_feat(287), I1 =>  inp_feat(242), I2 =>  inp_feat(183), I3 =>  inp_feat(448), I4 =>  inp_feat(77), I5 =>  inp_feat(402), I6 =>  inp_feat(29), I7 =>  inp_feat(58)); 
C_44_S_3_L_7_inst : LUT8 generic map(INIT => "0000110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001001101000000000000000000000000000001100000000000000000000000000100010000000000000001000000000000000000000000000000000000000000") port map( O =>C_44_S_3_L_7_out, I0 =>  inp_feat(457), I1 =>  inp_feat(407), I2 =>  inp_feat(204), I3 =>  inp_feat(237), I4 =>  inp_feat(259), I5 =>  inp_feat(477), I6 =>  inp_feat(296), I7 =>  inp_feat(384)); 
C_44_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000001000000100000000000100000000000001000000000000000000000000000001100101111000000001010101000000000000000000000000000110000000000000010000000100000101000100000000000000000000000000000000000000000101010000000000010101010") port map( O =>C_44_S_4_L_0_out, I0 =>  inp_feat(260), I1 =>  inp_feat(412), I2 =>  inp_feat(480), I3 =>  inp_feat(316), I4 =>  inp_feat(315), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_44_S_4_L_1_inst : LUT8 generic map(INIT => "1000001010100000111010001010000000000000000000000100000000000000000000000000101000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000") port map( O =>C_44_S_4_L_1_out, I0 =>  inp_feat(408), I1 =>  inp_feat(199), I2 =>  inp_feat(11), I3 =>  inp_feat(57), I4 =>  inp_feat(419), I5 =>  inp_feat(250), I6 =>  inp_feat(336), I7 =>  inp_feat(232)); 
C_44_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000001100010011001100010000000000101001001100110001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000") port map( O =>C_44_S_4_L_2_out, I0 =>  inp_feat(179), I1 =>  inp_feat(274), I2 =>  inp_feat(280), I3 =>  inp_feat(40), I4 =>  inp_feat(448), I5 =>  inp_feat(384), I6 =>  inp_feat(95), I7 =>  inp_feat(287)); 
C_44_S_4_L_3_inst : LUT8 generic map(INIT => "0000110000011000000111100000000000000000000000000000000001000000111010000011000011101100100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_4_L_3_out, I0 =>  inp_feat(334), I1 =>  inp_feat(504), I2 =>  inp_feat(432), I3 =>  inp_feat(180), I4 =>  inp_feat(73), I5 =>  inp_feat(34), I6 =>  inp_feat(452), I7 =>  inp_feat(183)); 
C_44_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000100000000000000000000000000000000000000000000000000111110100100000011101000100100001111000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_4_L_4_out, I0 =>  inp_feat(201), I1 =>  inp_feat(157), I2 =>  inp_feat(448), I3 =>  inp_feat(487), I4 =>  inp_feat(446), I5 =>  inp_feat(388), I6 =>  inp_feat(204), I7 =>  inp_feat(253)); 
C_44_S_4_L_5_inst : LUT8 generic map(INIT => "0000001011000110001000000111001100000000000000000000000001010101010100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_44_S_4_L_5_out, I0 =>  inp_feat(73), I1 =>  inp_feat(88), I2 =>  inp_feat(65), I3 =>  inp_feat(484), I4 =>  inp_feat(179), I5 =>  inp_feat(353), I6 =>  inp_feat(253), I7 =>  inp_feat(241)); 
C_44_S_4_L_6_inst : LUT8 generic map(INIT => "1000100010101000000000000000100000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000001000001000000000000010000000000000000000000000000000000000000000001000000000000000000000") port map( O =>C_44_S_4_L_6_out, I0 =>  inp_feat(487), I1 =>  inp_feat(171), I2 =>  inp_feat(162), I3 =>  inp_feat(92), I4 =>  inp_feat(362), I5 =>  inp_feat(347), I6 =>  inp_feat(172), I7 =>  inp_feat(459)); 
C_44_S_4_L_7_inst : LUT8 generic map(INIT => "0110000101111011000010001010101000000000000100010000000010000000000000001000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000") port map( O =>C_44_S_4_L_7_out, I0 =>  inp_feat(71), I1 =>  inp_feat(179), I2 =>  inp_feat(432), I3 =>  inp_feat(415), I4 =>  inp_feat(389), I5 =>  inp_feat(93), I6 =>  inp_feat(290), I7 =>  inp_feat(154)); 
C_45_S_0_L_0_inst : LUT8 generic map(INIT => "0010000000000000011000100011000100000000000000000010000000000000001010000000000010111010000000000000000000000000100000000000000000000000000000001010000000000000000000000000000000000000000000000010000000000000101100000000000000000000000000000000000000000000") port map( O =>C_45_S_0_L_0_out, I0 =>  inp_feat(322), I1 =>  inp_feat(445), I2 =>  inp_feat(407), I3 =>  inp_feat(153), I4 =>  inp_feat(316), I5 =>  inp_feat(487), I6 =>  inp_feat(419), I7 =>  inp_feat(2)); 
C_45_S_0_L_1_inst : LUT8 generic map(INIT => "0010000000000000101000000000000000000000000000000100000000000000111100000001000011110111011100010000000100000000011100110000000001110000011000001111100000000000100000000000000010000000000000001111000000000000101100000100000000000000000000000000000000000000") port map( O =>C_45_S_0_L_1_out, I0 =>  inp_feat(472), I1 =>  inp_feat(328), I2 =>  inp_feat(79), I3 =>  inp_feat(87), I4 =>  inp_feat(195), I5 =>  inp_feat(387), I6 =>  inp_feat(467), I7 =>  inp_feat(419)); 
C_45_S_0_L_2_inst : LUT8 generic map(INIT => "0010001001000010101000000000001010100000001000000010000000010000001000010000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_0_L_2_out, I0 =>  inp_feat(444), I1 =>  inp_feat(453), I2 =>  inp_feat(162), I3 =>  inp_feat(286), I4 =>  inp_feat(126), I5 =>  inp_feat(402), I6 =>  inp_feat(5), I7 =>  inp_feat(250)); 
C_45_S_0_L_3_inst : LUT8 generic map(INIT => "1101110000000101100000001000000011000000000000001110000000000000010110010001000000010000000000000000000000000000000000000000000000101100000000000000000000000000110100000000000000000000000000000011000100000001000000000000000000000000000000000000000000000000") port map( O =>C_45_S_0_L_3_out, I0 =>  inp_feat(52), I1 =>  inp_feat(509), I2 =>  inp_feat(402), I3 =>  inp_feat(486), I4 =>  inp_feat(336), I5 =>  inp_feat(128), I6 =>  inp_feat(420), I7 =>  inp_feat(286)); 
C_45_S_0_L_4_inst : LUT8 generic map(INIT => "0010000011000000010000001100000000000000110101000100000001000000000000010000000010000000000000000000000011000000010000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_45_S_0_L_4_out, I0 =>  inp_feat(109), I1 =>  inp_feat(387), I2 =>  inp_feat(206), I3 =>  inp_feat(53), I4 =>  inp_feat(50), I5 =>  inp_feat(247), I6 =>  inp_feat(6), I7 =>  inp_feat(123)); 
C_45_S_0_L_5_inst : LUT8 generic map(INIT => "1000110100000101100011010000000000000100000011010100100000000000000000000000000000000000000000001000000000000000000000000000000010000001100000001100010000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_0_L_5_out, I0 =>  inp_feat(109), I1 =>  inp_feat(206), I2 =>  inp_feat(221), I3 =>  inp_feat(353), I4 =>  inp_feat(475), I5 =>  inp_feat(6), I6 =>  inp_feat(123), I7 =>  inp_feat(5)); 
C_45_S_0_L_6_inst : LUT8 generic map(INIT => "1110010010000000010000001000000000000000000000000000000000000000010001001000000011000000110100000000000000000000000011000000000000000000000000000100000011000000010000000000000000000000000000000100010000000000110100000000000000000000000000000000000000000000") port map( O =>C_45_S_0_L_6_out, I0 =>  inp_feat(453), I1 =>  inp_feat(359), I2 =>  inp_feat(440), I3 =>  inp_feat(412), I4 =>  inp_feat(316), I5 =>  inp_feat(21), I6 =>  inp_feat(315), I7 =>  inp_feat(90)); 
C_45_S_0_L_7_inst : LUT8 generic map(INIT => "1000001010001010100000001000100010001000100010000000000010001000100010100000000000000010000000000100010011000101000000001000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000") port map( O =>C_45_S_0_L_7_out, I0 =>  inp_feat(130), I1 =>  inp_feat(357), I2 =>  inp_feat(411), I3 =>  inp_feat(73), I4 =>  inp_feat(397), I5 =>  inp_feat(247), I6 =>  inp_feat(6), I7 =>  inp_feat(123)); 
C_45_S_1_L_0_inst : LUT8 generic map(INIT => "0000100000000000000000100000000000000000000000000000000000000000001010110000000010001000000010000000101000000000000010000000100010101100000000000001100000001000000000000000000000001000100000001101111100000000100010000000100000001001000000000000101000000000") port map( O =>C_45_S_1_L_0_out, I0 =>  inp_feat(290), I1 =>  inp_feat(413), I2 =>  inp_feat(178), I3 =>  inp_feat(206), I4 =>  inp_feat(109), I5 =>  inp_feat(327), I6 =>  inp_feat(88), I7 =>  inp_feat(419)); 
C_45_S_1_L_1_inst : LUT8 generic map(INIT => "0011001000110000000000000101000000000000000100000000000000010000111110010111010000000000010100000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_1_L_1_out, I0 =>  inp_feat(329), I1 =>  inp_feat(317), I2 =>  inp_feat(387), I3 =>  inp_feat(380), I4 =>  inp_feat(87), I5 =>  inp_feat(416), I6 =>  inp_feat(61), I7 =>  inp_feat(250)); 
C_45_S_1_L_2_inst : LUT8 generic map(INIT => "0101101010110011010000000000000011101010000000100000001000000000100000100010101000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_1_L_2_out, I0 =>  inp_feat(134), I1 =>  inp_feat(88), I2 =>  inp_feat(272), I3 =>  inp_feat(109), I4 =>  inp_feat(5), I5 =>  inp_feat(232), I6 =>  inp_feat(59), I7 =>  inp_feat(250)); 
C_45_S_1_L_3_inst : LUT8 generic map(INIT => "0110100000100010100000000000000010101010001000100000000000000000000000000000100100000000000010000000001011101111000000000000101100001000000000000000000000000000000001000000010000000000000001000000000000001100000000000000100100000100000011000000010010101111") port map( O =>C_45_S_1_L_3_out, I0 =>  inp_feat(232), I1 =>  inp_feat(448), I2 =>  inp_feat(298), I3 =>  inp_feat(41), I4 =>  inp_feat(388), I5 =>  inp_feat(179), I6 =>  inp_feat(229), I7 =>  inp_feat(255)); 
C_45_S_1_L_4_inst : LUT8 generic map(INIT => "1001101010011010000001010000000100110010111100100010000000010000100000001000110000000000000000000000000010100000000000000000000000000000000000000000001000001000101000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_1_L_4_out, I0 =>  inp_feat(289), I1 =>  inp_feat(316), I2 =>  inp_feat(280), I3 =>  inp_feat(340), I4 =>  inp_feat(206), I5 =>  inp_feat(247), I6 =>  inp_feat(232), I7 =>  inp_feat(23)); 
C_45_S_1_L_5_inst : LUT8 generic map(INIT => "0000111000001100000000000000000010001110000000000000100000000000000000000000000000000100000000001000110000000000000000000000000010101010100000001010100000000000100111100100110010001010000000001000000000000000000000000000000000000100000001000000000000000000") port map( O =>C_45_S_1_L_5_out, I0 =>  inp_feat(420), I1 =>  inp_feat(29), I2 =>  inp_feat(316), I3 =>  inp_feat(86), I4 =>  inp_feat(164), I5 =>  inp_feat(247), I6 =>  inp_feat(23), I7 =>  inp_feat(340)); 
C_45_S_1_L_6_inst : LUT8 generic map(INIT => "0100000001000000000000001100000000000000110001100010000000000000010000000001011100100000000000010110001011010010001000000100000111000000110000000000000000000000110000101100000000100000000000000000000000000000000000000000000000100010100000000010001000000000") port map( O =>C_45_S_1_L_6_out, I0 =>  inp_feat(152), I1 =>  inp_feat(422), I2 =>  inp_feat(379), I3 =>  inp_feat(247), I4 =>  inp_feat(87), I5 =>  inp_feat(493), I6 =>  inp_feat(3), I7 =>  inp_feat(262)); 
C_45_S_1_L_7_inst : LUT8 generic map(INIT => "0000000010001000000100001110100010000001101101010001111011010100100100000101000011000000000100000000000000000000000000010100000000000000000010000000000000000000000000001000000101000001010100000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_1_L_7_out, I0 =>  inp_feat(130), I1 =>  inp_feat(251), I2 =>  inp_feat(342), I3 =>  inp_feat(221), I4 =>  inp_feat(36), I5 =>  inp_feat(403), I6 =>  inp_feat(87), I7 =>  inp_feat(66)); 
C_45_S_2_L_0_inst : LUT8 generic map(INIT => "1100100010000000110000000000000000000000000000001100000001000000111000001000000011000000100000000000000011000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_2_L_0_out, I0 =>  inp_feat(121), I1 =>  inp_feat(11), I2 =>  inp_feat(87), I3 =>  inp_feat(471), I4 =>  inp_feat(410), I5 =>  inp_feat(54), I6 =>  inp_feat(1), I7 =>  inp_feat(21)); 
C_45_S_2_L_1_inst : LUT8 generic map(INIT => "0100010001001000110011100010001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000011000001110011111000110000001100000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_2_L_1_out, I0 =>  inp_feat(472), I1 =>  inp_feat(132), I2 =>  inp_feat(378), I3 =>  inp_feat(6), I4 =>  inp_feat(55), I5 =>  inp_feat(42), I6 =>  inp_feat(250), I7 =>  inp_feat(479)); 
C_45_S_2_L_2_inst : LUT8 generic map(INIT => "0011000010100010000000000001000000100010101000000000000000001000110100001111000000010000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000") port map( O =>C_45_S_2_L_2_out, I0 =>  inp_feat(204), I1 =>  inp_feat(267), I2 =>  inp_feat(508), I3 =>  inp_feat(280), I4 =>  inp_feat(23), I5 =>  inp_feat(397), I6 =>  inp_feat(273), I7 =>  inp_feat(21)); 
C_45_S_2_L_3_inst : LUT8 generic map(INIT => "0101001010000000110010101000000011010100100000001000010010000000100000000000000011000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000") port map( O =>C_45_S_2_L_3_out, I0 =>  inp_feat(400), I1 =>  inp_feat(201), I2 =>  inp_feat(232), I3 =>  inp_feat(55), I4 =>  inp_feat(50), I5 =>  inp_feat(247), I6 =>  inp_feat(466), I7 =>  inp_feat(250)); 
C_45_S_2_L_4_inst : LUT8 generic map(INIT => "1101101001010111000000000100010100010101100101110000010100000101000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000001010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_2_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(340), I2 =>  inp_feat(419), I3 =>  inp_feat(448), I4 =>  inp_feat(45), I5 =>  inp_feat(247), I6 =>  inp_feat(232), I7 =>  inp_feat(23)); 
C_45_S_2_L_5_inst : LUT8 generic map(INIT => "0111101100001100000011001100110000000100100010000000001000000000000000000000000000000000000000000000000000000000000000000000000001101000100000010000011011001101000001000000110010001101000010010000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_45_S_2_L_5_out, I0 =>  inp_feat(445), I1 =>  inp_feat(170), I2 =>  inp_feat(448), I3 =>  inp_feat(73), I4 =>  inp_feat(179), I5 =>  inp_feat(229), I6 =>  inp_feat(192), I7 =>  inp_feat(298)); 
C_45_S_2_L_6_inst : LUT8 generic map(INIT => "0000100010000000011000100000000001000000000000000000000000000000010011010100000000000000000000001000000000000000000000000000000000000000100000001011101000000000110000000000000000000000000000001100000010000000000000000000100000000000000000000000100000001000") port map( O =>C_45_S_2_L_6_out, I0 =>  inp_feat(420), I1 =>  inp_feat(407), I2 =>  inp_feat(354), I3 =>  inp_feat(73), I4 =>  inp_feat(451), I5 =>  inp_feat(287), I6 =>  inp_feat(64), I7 =>  inp_feat(1)); 
C_45_S_2_L_7_inst : LUT8 generic map(INIT => "0010100000001010111010100000101010000000100010000000000010001010000000000000000000000000101110000000000010001000000000101100110000000000001000000000000010110000100000001010000000000000110001000000000000000000000000001100010000000000000000000000000001000100") port map( O =>C_45_S_2_L_7_out, I0 =>  inp_feat(388), I1 =>  inp_feat(103), I2 =>  inp_feat(267), I3 =>  inp_feat(317), I4 =>  inp_feat(404), I5 =>  inp_feat(340), I6 =>  inp_feat(229), I7 =>  inp_feat(76)); 
C_45_S_3_L_0_inst : LUT8 generic map(INIT => "1110001100000000100011000000100010000001000000011000000000000000000000100000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000") port map( O =>C_45_S_3_L_0_out, I0 =>  inp_feat(460), I1 =>  inp_feat(400), I2 =>  inp_feat(247), I3 =>  inp_feat(503), I4 =>  inp_feat(131), I5 =>  inp_feat(232), I6 =>  inp_feat(23), I7 =>  inp_feat(250)); 
C_45_S_3_L_1_inst : LUT8 generic map(INIT => "0111000000100000000000000000000000000000010000000000000000000000101100111010101100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_3_L_1_out, I0 =>  inp_feat(374), I1 =>  inp_feat(40), I2 =>  inp_feat(426), I3 =>  inp_feat(11), I4 =>  inp_feat(232), I5 =>  inp_feat(359), I6 =>  inp_feat(55), I7 =>  inp_feat(21)); 
C_45_S_3_L_2_inst : LUT8 generic map(INIT => "0111011010010100000000000100000001110010001000000010000000000000011100001100000100000000000000000111100100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000") port map( O =>C_45_S_3_L_2_out, I0 =>  inp_feat(472), I1 =>  inp_feat(317), I2 =>  inp_feat(87), I3 =>  inp_feat(475), I4 =>  inp_feat(83), I5 =>  inp_feat(232), I6 =>  inp_feat(473), I7 =>  inp_feat(21)); 
C_45_S_3_L_3_inst : LUT8 generic map(INIT => "1111111101110001000000000000000000010000000000000000000000000000101100110000000000000010000000000000010000000000000000000000000001110101100000000000000000000000000000000000000000000000000000000011010100010100000000000000000000001100000000000000000000000000") port map( O =>C_45_S_3_L_3_out, I0 =>  inp_feat(340), I1 =>  inp_feat(1), I2 =>  inp_feat(336), I3 =>  inp_feat(251), I4 =>  inp_feat(42), I5 =>  inp_feat(209), I6 =>  inp_feat(298), I7 =>  inp_feat(364)); 
C_45_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000010001000100010011000000000000000000000000000000000000000100000010100100100000110100010000000000000000000010000000000001110000000000000001000001010000000000000000000000000000000000000101100010000000010110000001000000001000000000000000100000000000") port map( O =>C_45_S_3_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(316), I2 =>  inp_feat(336), I3 =>  inp_feat(74), I4 =>  inp_feat(109), I5 =>  inp_feat(188), I6 =>  inp_feat(41), I7 =>  inp_feat(262)); 
C_45_S_3_L_5_inst : LUT8 generic map(INIT => "0100000000001100100001100100010000011100110000001010110101001100001000000000000000000000000001000000000000000000000011010000100000000000010100010000000000000000000010000000000000001000000000000000000000000001100010111000111100000000000000000000100000001000") port map( O =>C_45_S_3_L_5_out, I0 =>  inp_feat(461), I1 =>  inp_feat(85), I2 =>  inp_feat(115), I3 =>  inp_feat(109), I4 =>  inp_feat(311), I5 =>  inp_feat(430), I6 =>  inp_feat(192), I7 =>  inp_feat(255)); 
C_45_S_3_L_6_inst : LUT8 generic map(INIT => "1010000000100000000000000000000000000000000000000000000000000000101100001110000000000000000000000000000000000000000000000000000000100010111000100000000011100000000000000000000000000000000000001011000001010001111000001101000010000000000100010100000000000000") port map( O =>C_45_S_3_L_6_out, I0 =>  inp_feat(488), I1 =>  inp_feat(115), I2 =>  inp_feat(482), I3 =>  inp_feat(85), I4 =>  inp_feat(155), I5 =>  inp_feat(306), I6 =>  inp_feat(30), I7 =>  inp_feat(417)); 
C_45_S_3_L_7_inst : LUT8 generic map(INIT => "0010000010110011111000000000000001000000000000000000000001001100000000001000100000000000000000000000000010000010000000000000000010110101001101010100000100010101010000000000000000000000110011000000000000001001000101000001111000100010001000100000100000001100") port map( O =>C_45_S_3_L_7_out, I0 =>  inp_feat(298), I1 =>  inp_feat(461), I2 =>  inp_feat(11), I3 =>  inp_feat(430), I4 =>  inp_feat(93), I5 =>  inp_feat(449), I6 =>  inp_feat(34), I7 =>  inp_feat(266)); 
C_45_S_4_L_0_inst : LUT8 generic map(INIT => "0000000100000000000100000000000011010000100000000001000000010000000000000000000000000000000000000000100000001000000000000000000011100000000000000001000000000000111000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_45_S_4_L_0_out, I0 =>  inp_feat(374), I1 =>  inp_feat(152), I2 =>  inp_feat(344), I3 =>  inp_feat(206), I4 =>  inp_feat(160), I5 =>  inp_feat(109), I6 =>  inp_feat(250), I7 =>  inp_feat(328)); 
C_45_S_4_L_1_inst : LUT8 generic map(INIT => "0100100000000000111000000000000001000001000000000000000000000000100000001000000001000000000000000000111000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010") port map( O =>C_45_S_4_L_1_out, I0 =>  inp_feat(176), I1 =>  inp_feat(23), I2 =>  inp_feat(45), I3 =>  inp_feat(286), I4 =>  inp_feat(229), I5 =>  inp_feat(131), I6 =>  inp_feat(109), I7 =>  inp_feat(250)); 
C_45_S_4_L_2_inst : LUT8 generic map(INIT => "1100000110000000100110011000000000001101000000001000000010000000000000001000000011011001100000000000000000000000000000001000000010000010000000000011000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000") port map( O =>C_45_S_4_L_2_out, I0 =>  inp_feat(186), I1 =>  inp_feat(403), I2 =>  inp_feat(172), I3 =>  inp_feat(131), I4 =>  inp_feat(448), I5 =>  inp_feat(54), I6 =>  inp_feat(87), I7 =>  inp_feat(387)); 
C_45_S_4_L_3_inst : LUT8 generic map(INIT => "0000100000000100000000000000000001010011000000000000000000000000011100110100000001010000000000000011001100000000001000011000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000") port map( O =>C_45_S_4_L_3_out, I0 =>  inp_feat(480), I1 =>  inp_feat(30), I2 =>  inp_feat(20), I3 =>  inp_feat(344), I4 =>  inp_feat(206), I5 =>  inp_feat(160), I6 =>  inp_feat(109), I7 =>  inp_feat(250)); 
C_45_S_4_L_4_inst : LUT8 generic map(INIT => "0110010001101110011000000000011000000000000010001000000000001000011010000001100010000000000000001110000011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_45_S_4_L_4_out, I0 =>  inp_feat(380), I1 =>  inp_feat(14), I2 =>  inp_feat(6), I3 =>  inp_feat(378), I4 =>  inp_feat(85), I5 =>  inp_feat(131), I6 =>  inp_feat(109), I7 =>  inp_feat(250)); 
C_45_S_4_L_5_inst : LUT8 generic map(INIT => "1100110001001100000010000000000000000101000000000000100000001000110011010000100000000000110010000000010100000000000000000000000011111101110011000000000000000000100001000000000000000000000000000111010100000000000000001000100001010101000000000000000000000000") port map( O =>C_45_S_4_L_5_out, I0 =>  inp_feat(266), I1 =>  inp_feat(87), I2 =>  inp_feat(262), I3 =>  inp_feat(410), I4 =>  inp_feat(157), I5 =>  inp_feat(271), I6 =>  inp_feat(252), I7 =>  inp_feat(198)); 
C_45_S_4_L_6_inst : LUT8 generic map(INIT => "1100110000000000100000001000000001000000000000000000000000000000010011000010000110000101000001010000000000000000000000000000000001001001000000000000000000000000000000000000000000100000000000000110110110001011000010101000110100000000000000000000000000000000") port map( O =>C_45_S_4_L_6_out, I0 =>  inp_feat(267), I1 =>  inp_feat(232), I2 =>  inp_feat(493), I3 =>  inp_feat(166), I4 =>  inp_feat(477), I5 =>  inp_feat(95), I6 =>  inp_feat(479), I7 =>  inp_feat(198)); 
C_45_S_4_L_7_inst : LUT8 generic map(INIT => "1101000000010000110100000001000001000000000000000111000000000000100010001000000010000000000000001000100000000000000100000000000010000010000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000") port map( O =>C_45_S_4_L_7_out, I0 =>  inp_feat(73), I1 =>  inp_feat(301), I2 =>  inp_feat(388), I3 =>  inp_feat(35), I4 =>  inp_feat(365), I5 =>  inp_feat(229), I6 =>  inp_feat(19), I7 =>  inp_feat(5)); 
C_46_S_0_L_0_inst : LUT8 generic map(INIT => "1111111111101010111101011111111101110010010000001101000001010000001110101000100001000000111000000000000000000000000000000100000000000000100000001100000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_46_S_0_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(265), I2 =>  inp_feat(317), I3 =>  inp_feat(496), I4 =>  inp_feat(27), I5 =>  inp_feat(484), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_46_S_0_L_1_inst : LUT8 generic map(INIT => "1110001011111011000000001110100011000010000000000000000010000000111000101010101010000000101000001110001000000000000000001000000011110000111101110011000001111010011101100000000000000000000000000010000000000000000000000000000011111010000000000000000000000000") port map( O =>C_46_S_0_L_1_out, I0 =>  inp_feat(37), I1 =>  inp_feat(302), I2 =>  inp_feat(134), I3 =>  inp_feat(336), I4 =>  inp_feat(419), I5 =>  inp_feat(253), I6 =>  inp_feat(388), I7 =>  inp_feat(211)); 
C_46_S_0_L_2_inst : LUT8 generic map(INIT => "1110101011001010101010100000100011101111101010100000101000001010000001000000100000000010000000001010101100001000000010000000100011111111000010001010101000000000101111110000101000000000000000001001111100000000000000000000000010011111000000000000000000000000") port map( O =>C_46_S_0_L_2_out, I0 =>  inp_feat(258), I1 =>  inp_feat(383), I2 =>  inp_feat(494), I3 =>  inp_feat(485), I4 =>  inp_feat(284), I5 =>  inp_feat(171), I6 =>  inp_feat(484), I7 =>  inp_feat(183)); 
C_46_S_0_L_3_inst : LUT8 generic map(INIT => "1111111001110100111110101111000011010000010100001000000011000000001011000000000000000000100000000000000011000000000000000000000011111100111101111111100011001000000000000010000011000000110000000100110010000000100000001100000000000000010000001100000011000000") port map( O =>C_46_S_0_L_3_out, I0 =>  inp_feat(201), I1 =>  inp_feat(51), I2 =>  inp_feat(183), I3 =>  inp_feat(75), I4 =>  inp_feat(130), I5 =>  inp_feat(276), I6 =>  inp_feat(235), I7 =>  inp_feat(302)); 
C_46_S_0_L_4_inst : LUT8 generic map(INIT => "1010011010110000101011001010000011111110010100000000111000000000101010100001000000100010000000001011101000010000000000000000000000100010000000001000001010000000101000100000000000000010000000001010100000010000101000100000000000110010001100000010001000000000") port map( O =>C_46_S_0_L_4_out, I0 =>  inp_feat(415), I1 =>  inp_feat(427), I2 =>  inp_feat(411), I3 =>  inp_feat(126), I4 =>  inp_feat(379), I5 =>  inp_feat(302), I6 =>  inp_feat(264), I7 =>  inp_feat(273)); 
C_46_S_0_L_5_inst : LUT8 generic map(INIT => "1000101010000000000000001000000010001000100000001000101010000000101000011000000000001010000000001010000010000000000010100000000010101010001010000000100000000000101010100000000000001010000000000000001000000000000010100000000010001010000000000000101000000000") port map( O =>C_46_S_0_L_5_out, I0 =>  inp_feat(2), I1 =>  inp_feat(204), I2 =>  inp_feat(270), I3 =>  inp_feat(284), I4 =>  inp_feat(63), I5 =>  inp_feat(435), I6 =>  inp_feat(296), I7 =>  inp_feat(444)); 
C_46_S_0_L_6_inst : LUT8 generic map(INIT => "0010110010000100101010101010101000001000100010001010100010101010110000001110111111001100000010000000000000001000100000000000000010001100101011100000101000001010000000000000000000000000000000001010100010101010100010000000100010000000000000000000000000000000") port map( O =>C_46_S_0_L_6_out, I0 =>  inp_feat(263), I1 =>  inp_feat(402), I2 =>  inp_feat(201), I3 =>  inp_feat(330), I4 =>  inp_feat(289), I5 =>  inp_feat(284), I6 =>  inp_feat(444), I7 =>  inp_feat(407)); 
C_46_S_0_L_7_inst : LUT8 generic map(INIT => "1111000001100100111000001111000010000000111011001010000010110000110001000100110011000000110111010000000000000000000000000000000011100000001000001000000000100000000000001000000000000000100000001100100011000001100000001100100000000000100000000000000000000000") port map( O =>C_46_S_0_L_7_out, I0 =>  inp_feat(88), I1 =>  inp_feat(225), I2 =>  inp_feat(366), I3 =>  inp_feat(201), I4 =>  inp_feat(108), I5 =>  inp_feat(244), I6 =>  inp_feat(183), I7 =>  inp_feat(384)); 
C_46_S_1_L_0_inst : LUT8 generic map(INIT => "1111111111101010111101011111111101110010010000001101000001010000001110101000100001000000111000000000000000000000000000000100000000000000100000001100000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_46_S_1_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(265), I2 =>  inp_feat(317), I3 =>  inp_feat(496), I4 =>  inp_feat(27), I5 =>  inp_feat(484), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_46_S_1_L_1_inst : LUT8 generic map(INIT => "1111100010100000111110001000000011100000101000001111000010100000111100010000000010110000100000001010000000100000100000000000000010000000000000001000100000000000110011011000000110000000101000000000000000000000101000000000000010000000100000001000000000100000") port map( O =>C_46_S_1_L_1_out, I0 =>  inp_feat(288), I1 =>  inp_feat(115), I2 =>  inp_feat(235), I3 =>  inp_feat(1), I4 =>  inp_feat(87), I5 =>  inp_feat(172), I6 =>  inp_feat(74), I7 =>  inp_feat(211)); 
C_46_S_1_L_2_inst : LUT8 generic map(INIT => "0101100011111000000110000000101010011100100011000000000000000100111110001111000010001000101000001101110000000000000000000000000011011000100000001000100010001000000110000000100000000000000000001101000000000000000010001000100001011100000000000000000000000000") port map( O =>C_46_S_1_L_2_out, I0 =>  inp_feat(350), I1 =>  inp_feat(284), I2 =>  inp_feat(444), I3 =>  inp_feat(387), I4 =>  inp_feat(320), I5 =>  inp_feat(336), I6 =>  inp_feat(34), I7 =>  inp_feat(183)); 
C_46_S_1_L_3_inst : LUT8 generic map(INIT => "0100100010100010001000001010101010001000100000001000000000000000111111001010000010000000000000001000000010100000000000000000000011101110000000001010100010101000100010000000000010000000000000001111000000000000000000000000000000000000000000000000000000000000") port map( O =>C_46_S_1_L_3_out, I0 =>  inp_feat(179), I1 =>  inp_feat(53), I2 =>  inp_feat(230), I3 =>  inp_feat(487), I4 =>  inp_feat(320), I5 =>  inp_feat(68), I6 =>  inp_feat(232), I7 =>  inp_feat(302)); 
C_46_S_1_L_4_inst : LUT8 generic map(INIT => "1100101011110000000000100010000011101100101000001010101010101010101000001100000010000010000000001010101000000000101010100010001000000000111000000000000000000000000010001010000010000010000000000000000011100000000000101000000000000000100000001010101010001000") port map( O =>C_46_S_1_L_4_out, I0 =>  inp_feat(504), I1 =>  inp_feat(484), I2 =>  inp_feat(383), I3 =>  inp_feat(27), I4 =>  inp_feat(320), I5 =>  inp_feat(302), I6 =>  inp_feat(264), I7 =>  inp_feat(273)); 
C_46_S_1_L_5_inst : LUT8 generic map(INIT => "1011101110001000001100010000100011111000100010000000000000000000101010100000100000000000000010001110100000001000101010000000000000110000000010000001000000000000111010000000100000001000100010001011101000001000000000000000100010001000000010001000100000001000") port map( O =>C_46_S_1_L_5_out, I0 =>  inp_feat(419), I1 =>  inp_feat(51), I2 =>  inp_feat(120), I3 =>  inp_feat(17), I4 =>  inp_feat(50), I5 =>  inp_feat(264), I6 =>  inp_feat(446), I7 =>  inp_feat(92)); 
C_46_S_1_L_6_inst : LUT8 generic map(INIT => "1010001010110000111100001111000011110011100000001001001110000000101000110001000010110001001100001000100000000000100010110000000000100010000000000000000000000000001100101000000000010000000000000000000000000010000100000000000000100000000000000000000100000000") port map( O =>C_46_S_1_L_6_out, I0 =>  inp_feat(445), I1 =>  inp_feat(494), I2 =>  inp_feat(415), I3 =>  inp_feat(73), I4 =>  inp_feat(264), I5 =>  inp_feat(331), I6 =>  inp_feat(134), I7 =>  inp_feat(425)); 
C_46_S_1_L_7_inst : LUT8 generic map(INIT => "1101010010001010110110001000000011010000110000001111001000000000111111010000000011101101000000000000000000000000101010000000000011111010101010101000101000000010111110101110101001101010101010101100111000000000110000000000000010100010000000000000000000000000") port map( O =>C_46_S_1_L_7_out, I0 =>  inp_feat(130), I1 =>  inp_feat(484), I2 =>  inp_feat(151), I3 =>  inp_feat(442), I4 =>  inp_feat(157), I5 =>  inp_feat(5), I6 =>  inp_feat(34), I7 =>  inp_feat(183)); 
C_46_S_2_L_0_inst : LUT8 generic map(INIT => "1111111111101010111101011111111101110010010000001101000001010000001110101000100001000000111000000000000000000000000000000100000000000000100000001100000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_46_S_2_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(265), I2 =>  inp_feat(317), I3 =>  inp_feat(496), I4 =>  inp_feat(27), I5 =>  inp_feat(484), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_46_S_2_L_1_inst : LUT8 generic map(INIT => "1111111110100010101000001010001011110100001000001010000000100010101010000000000010000000000000101000100000000000000000000000001011111110000000001011000010000000110000000000000000000000000000001110111100000000101100001000000011000000000000000000000000000000") port map( O =>C_46_S_2_L_1_out, I0 =>  inp_feat(204), I1 =>  inp_feat(178), I2 =>  inp_feat(448), I3 =>  inp_feat(315), I4 =>  inp_feat(68), I5 =>  inp_feat(20), I6 =>  inp_feat(484), I7 =>  inp_feat(287)); 
C_46_S_2_L_2_inst : LUT8 generic map(INIT => "1111111100001100000001000000000011001111010001001000010100000000101111111100110010001111100011001000111100000000000000110000000010001101100010001000000000000000100000000000000011000000000000001000110010000000000010100000000000000110000000000000001100000000") port map( O =>C_46_S_2_L_2_out, I0 =>  inp_feat(142), I1 =>  inp_feat(187), I2 =>  inp_feat(171), I3 =>  inp_feat(134), I4 =>  inp_feat(109), I5 =>  inp_feat(259), I6 =>  inp_feat(172), I7 =>  inp_feat(183)); 
C_46_S_2_L_3_inst : LUT8 generic map(INIT => "0000001011001010101100001000100010111011100010111011000010000000101010101000101000000000100000001010101000001011000000000000000010110010010000100101000000000000001110111000100001010000000000001010101000100010000000000000000010100010101000100000000000000000") port map( O =>C_46_S_2_L_3_out, I0 =>  inp_feat(262), I1 =>  inp_feat(302), I2 =>  inp_feat(245), I3 =>  inp_feat(379), I4 =>  inp_feat(487), I5 =>  inp_feat(387), I6 =>  inp_feat(172), I7 =>  inp_feat(12)); 
C_46_S_2_L_4_inst : LUT8 generic map(INIT => "1110111011101011101110110001111100101010101000001000000000000000000011111010111100000000000000001000110010000000000000000000000011001110100000000000010000000000110111110000000000000000000000001100110000000000000000000000000011111111000000000000000000000000") port map( O =>C_46_S_2_L_4_out, I0 =>  inp_feat(109), I1 =>  inp_feat(26), I2 =>  inp_feat(71), I3 =>  inp_feat(379), I4 =>  inp_feat(284), I5 =>  inp_feat(406), I6 =>  inp_feat(331), I7 =>  inp_feat(354)); 
C_46_S_2_L_5_inst : LUT8 generic map(INIT => "0111111100100100111011011010111111110000000000001111000000000000000111110000000000000001000000001000000000000000000000000000000010101111000001111010111100101111101000000000000010100010000000000000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_46_S_2_L_5_out, I0 =>  inp_feat(274), I1 =>  inp_feat(201), I2 =>  inp_feat(456), I3 =>  inp_feat(490), I4 =>  inp_feat(444), I5 =>  inp_feat(51), I6 =>  inp_feat(284), I7 =>  inp_feat(446)); 
C_46_S_2_L_6_inst : LUT8 generic map(INIT => "1111111111100100110011010100000000000111000000000000000000000000000101010000000000000000000000000101010100000000000000000000000010101111100010000010100100000000100000010000000000000000000000000000000110001000000000000000000001110111000000000000000000000000") port map( O =>C_46_S_2_L_6_out, I0 =>  inp_feat(302), I1 =>  inp_feat(75), I2 =>  inp_feat(509), I3 =>  inp_feat(50), I4 =>  inp_feat(273), I5 =>  inp_feat(18), I6 =>  inp_feat(299), I7 =>  inp_feat(229)); 
C_46_S_2_L_7_inst : LUT8 generic map(INIT => "0000110010101010000000001000110010001110101010100000011010001000100000001000101000000000000010101000000010000000100000001010101011100010111000110000000000001100000011100000101100001110100010000000000010101010000000000000000000000000001000110000000010101011") port map( O =>C_46_S_2_L_7_out, I0 =>  inp_feat(425), I1 =>  inp_feat(273), I2 =>  inp_feat(494), I3 =>  inp_feat(7), I4 =>  inp_feat(384), I5 =>  inp_feat(302), I6 =>  inp_feat(264), I7 =>  inp_feat(274)); 
C_46_S_3_L_0_inst : LUT8 generic map(INIT => "1111111111101010111101011111111101110010010000001101000001010000001110101000100001000000111000000000000000000000000000000100000000000000100000001100000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_46_S_3_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(265), I2 =>  inp_feat(317), I3 =>  inp_feat(496), I4 =>  inp_feat(27), I5 =>  inp_feat(484), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_46_S_3_L_1_inst : LUT8 generic map(INIT => "1000100000000000101010101000000011111011101010001010111010000000110000001000000010000000000000001110000010000000101010100000000011101100100000001000000000000000001100001000000010000010100000001100000000000000100000000000000000000000000000001000000000000000") port map( O =>C_46_S_3_L_1_out, I0 =>  inp_feat(366), I1 =>  inp_feat(152), I2 =>  inp_feat(504), I3 =>  inp_feat(134), I4 =>  inp_feat(172), I5 =>  inp_feat(336), I6 =>  inp_feat(132), I7 =>  inp_feat(287)); 
C_46_S_3_L_2_inst : LUT8 generic map(INIT => "1011111110111011101010101010001000000000001100001010000010100000100010011010000110000000100000000000000011000000000000001000000010111011101100111010001010101010100000000001000000000000000000001001011111110111100000001000000000000000110000000000000010000000") port map( O =>C_46_S_3_L_2_out, I0 =>  inp_feat(92), I1 =>  inp_feat(302), I2 =>  inp_feat(264), I3 =>  inp_feat(154), I4 =>  inp_feat(34), I5 =>  inp_feat(178), I6 =>  inp_feat(50), I7 =>  inp_feat(183)); 
C_46_S_3_L_3_inst : LUT8 generic map(INIT => "1111101011100010110000000000000011101010000000001000100000000000101010100010000000000000000000001010101000000000100010000000000011101010010000000100000001000000110000001000000011000000010000000010001010000000000000000000000000001000000000000000000000000000") port map( O =>C_46_S_3_L_3_out, I0 =>  inp_feat(288), I1 =>  inp_feat(27), I2 =>  inp_feat(452), I3 =>  inp_feat(412), I4 =>  inp_feat(50), I5 =>  inp_feat(183), I6 =>  inp_feat(316), I7 =>  inp_feat(419)); 
C_46_S_3_L_4_inst : LUT8 generic map(INIT => "1111100001101010011000100010101010100100111000000000000000000000101100101110101011100000111010100010000011100000001000000000000000001100001000000000000000000000000000000000000000000000000000001010000000100010101000000000000000100000001000000010000000000000") port map( O =>C_46_S_3_L_4_out, I0 =>  inp_feat(504), I1 =>  inp_feat(302), I2 =>  inp_feat(179), I3 =>  inp_feat(130), I4 =>  inp_feat(452), I5 =>  inp_feat(397), I6 =>  inp_feat(406), I7 =>  inp_feat(214)); 
C_46_S_3_L_5_inst : LUT8 generic map(INIT => "1010100010001110101011100000100110100000111010101000010000000010100011111000111000000000000011001000011011001111000000000000111111001100110011000000100000000000000000001100000000000000000000000000000000000000000000000000000010000000110000000000000000000000") port map( O =>C_46_S_3_L_5_out, I0 =>  inp_feat(484), I1 =>  inp_feat(412), I2 =>  inp_feat(494), I3 =>  inp_feat(171), I4 =>  inp_feat(179), I5 =>  inp_feat(406), I6 =>  inp_feat(411), I7 =>  inp_feat(423)); 
C_46_S_3_L_6_inst : LUT8 generic map(INIT => "1010000011110000111101000100000010000000101000001001000010100000111001000000000001000100000000001110010010000000111000001010000011001100110001000000000000000000111001000000000000100000101000000100000000000000000000000000000011000100001000001110010010100000") port map( O =>C_46_S_3_L_6_out, I0 =>  inp_feat(221), I1 =>  inp_feat(204), I2 =>  inp_feat(315), I3 =>  inp_feat(264), I4 =>  inp_feat(383), I5 =>  inp_feat(456), I6 =>  inp_feat(253), I7 =>  inp_feat(97)); 
C_46_S_3_L_7_inst : LUT8 generic map(INIT => "1111001011111100100000001010000011000000101010001000000000000000000000000000000000000000000000001100000000000000000010000000100011111010111011101100100000001000111010001010100011001000000010000000100000101000000000000000100010001000101010000000100000001000") port map( O =>C_46_S_3_L_7_out, I0 =>  inp_feat(88), I1 =>  inp_feat(411), I2 =>  inp_feat(134), I3 =>  inp_feat(264), I4 =>  inp_feat(92), I5 =>  inp_feat(183), I6 =>  inp_feat(490), I7 =>  inp_feat(302)); 
C_46_S_4_L_0_inst : LUT8 generic map(INIT => "1111111111101010111101011111111101110010010000001101000001010000001110101000100001000000111000000000000000000000000000000100000000000000100000001100000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_46_S_4_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(265), I2 =>  inp_feat(317), I3 =>  inp_feat(496), I4 =>  inp_feat(27), I5 =>  inp_feat(484), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_46_S_4_L_1_inst : LUT8 generic map(INIT => "1000100000000000101010101000000011111011101010001010111010000000110000001000000010000000000000001110000010000000101010100000000011101100100000001000000000000000001100001000000010000010100000001100000000000000100000000000000000000000000000001000000000000000") port map( O =>C_46_S_4_L_1_out, I0 =>  inp_feat(366), I1 =>  inp_feat(152), I2 =>  inp_feat(504), I3 =>  inp_feat(134), I4 =>  inp_feat(172), I5 =>  inp_feat(336), I6 =>  inp_feat(132), I7 =>  inp_feat(287)); 
C_46_S_4_L_2_inst : LUT8 generic map(INIT => "1011111110111011101010101010001000000000001100001010000010100000100010011010000110000000100000000000000011000000000000001000000010111011101100111010001010101010100000000001000000000000000000001001011111110111100000001000000000000000110000000000000010000000") port map( O =>C_46_S_4_L_2_out, I0 =>  inp_feat(92), I1 =>  inp_feat(302), I2 =>  inp_feat(264), I3 =>  inp_feat(154), I4 =>  inp_feat(34), I5 =>  inp_feat(178), I6 =>  inp_feat(50), I7 =>  inp_feat(183)); 
C_46_S_4_L_3_inst : LUT8 generic map(INIT => "1111101101110001101110110000001010111010001100001011101000111010111100000010100000111010001100101011000011110000101110101011101010100000000000100000101000000000100000100000000010100010001000101000000000000000000010100000000000000000000000000000000000100000") port map( O =>C_46_S_4_L_3_out, I0 =>  inp_feat(402), I1 =>  inp_feat(302), I2 =>  inp_feat(212), I3 =>  inp_feat(484), I4 =>  inp_feat(171), I5 =>  inp_feat(438), I6 =>  inp_feat(452), I7 =>  inp_feat(419)); 
C_46_S_4_L_4_inst : LUT8 generic map(INIT => "0010011100101111101001101010001010011000001000010000000000100000010110111010011111001100101000000111111110100011000000001010000001110100100011000000000010101000011111001110110000000000000000001000000010000000000000000000000000000000001000000000000000000000") port map( O =>C_46_S_4_L_4_out, I0 =>  inp_feat(37), I1 =>  inp_feat(407), I2 =>  inp_feat(334), I3 =>  inp_feat(302), I4 =>  inp_feat(314), I5 =>  inp_feat(242), I6 =>  inp_feat(264), I7 =>  inp_feat(54)); 
C_46_S_4_L_5_inst : LUT8 generic map(INIT => "1110110010001000000000001000100011101010100010000000000010001000111101011000000000010010100000001111111110000000100000001000000011101110110011001010000010000000100000101000100000001000100010001000010010000000100000001000000010000000100000001010000010001000") port map( O =>C_46_S_4_L_5_out, I0 =>  inp_feat(119), I1 =>  inp_feat(334), I2 =>  inp_feat(383), I3 =>  inp_feat(183), I4 =>  inp_feat(484), I5 =>  inp_feat(388), I6 =>  inp_feat(54), I7 =>  inp_feat(5)); 
C_46_S_4_L_6_inst : LUT8 generic map(INIT => "1010000011011100111110000001100011011000111000001110000000000000111010001110000010110000000000001110000011110000000000000000000011001100010111001111110011101000101000001100000010100000100000001000000011000000001000001010000011000000111100000000000000000000") port map( O =>C_46_S_4_L_6_out, I0 =>  inp_feat(484), I1 =>  inp_feat(273), I2 =>  inp_feat(169), I3 =>  inp_feat(134), I4 =>  inp_feat(346), I5 =>  inp_feat(331), I6 =>  inp_feat(264), I7 =>  inp_feat(97)); 
C_46_S_4_L_7_inst : LUT8 generic map(INIT => "1100110101010001011110001011000011000100000000000000000010100000111011010011011110101000101000001000110000000000000000000010000000000000010000010100000001000000000000000000000000100000000000001000110001000101000000000110000000000000000000000000000000000000") port map( O =>C_46_S_4_L_7_out, I0 =>  inp_feat(427), I1 =>  inp_feat(450), I2 =>  inp_feat(298), I3 =>  inp_feat(242), I4 =>  inp_feat(54), I5 =>  inp_feat(14), I6 =>  inp_feat(302), I7 =>  inp_feat(320)); 
C_47_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000001111111010001000000000000000000000000000000010000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000100010000000000000000000") port map( O =>C_47_S_0_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(373), I2 =>  inp_feat(355), I3 =>  inp_feat(82), I4 =>  inp_feat(34), I5 =>  inp_feat(221), I6 =>  inp_feat(199), I7 =>  inp_feat(2)); 
C_47_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111011000110110000000000100000000000000000000000000010000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_0_L_1_out, I0 =>  inp_feat(99), I1 =>  inp_feat(408), I2 =>  inp_feat(307), I3 =>  inp_feat(93), I4 =>  inp_feat(476), I5 =>  inp_feat(338), I6 =>  inp_feat(251), I7 =>  inp_feat(345)); 
C_47_S_0_L_2_inst : LUT8 generic map(INIT => "0000000100000100000000000000000000001100000001010000100000000000110110100000000011100000000000000000111100001101000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000110000000000000000000") port map( O =>C_47_S_0_L_2_out, I0 =>  inp_feat(301), I1 =>  inp_feat(161), I2 =>  inp_feat(221), I3 =>  inp_feat(365), I4 =>  inp_feat(387), I5 =>  inp_feat(448), I6 =>  inp_feat(452), I7 =>  inp_feat(87)); 
C_47_S_0_L_3_inst : LUT8 generic map(INIT => "0000000100000000001000010000000000100010100000000010001100000000000000000000000000000010000000000000000000000000000100110000000010100000000100001010000000000000101000000111000000100010000000000000000000000000001000000000000000000000000000000000000000000000") port map( O =>C_47_S_0_L_3_out, I0 =>  inp_feat(84), I1 =>  inp_feat(380), I2 =>  inp_feat(158), I3 =>  inp_feat(128), I4 =>  inp_feat(36), I5 =>  inp_feat(504), I6 =>  inp_feat(100), I7 =>  inp_feat(419)); 
C_47_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000110000000000001001000011001000000100000000000010100011000000000000000000000000000000000000000000000000000000001000000010000000101110101010100000100000000000001010000010100000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_0_L_4_out, I0 =>  inp_feat(407), I1 =>  inp_feat(92), I2 =>  inp_feat(154), I3 =>  inp_feat(316), I4 =>  inp_feat(178), I5 =>  inp_feat(419), I6 =>  inp_feat(287), I7 =>  inp_feat(134)); 
C_47_S_0_L_5_inst : LUT8 generic map(INIT => "1011001000000000001000000000000000000000001000000000000000000000001000000000000000000000000000000000001000000000000000000000000010110010100000000010101000000000001100000010000000010000000000000000001000000000001000100000000000110000000000000000000000000000") port map( O =>C_47_S_0_L_5_out, I0 =>  inp_feat(424), I1 =>  inp_feat(384), I2 =>  inp_feat(387), I3 =>  inp_feat(407), I4 =>  inp_feat(296), I5 =>  inp_feat(354), I6 =>  inp_feat(388), I7 =>  inp_feat(445)); 
C_47_S_0_L_6_inst : LUT8 generic map(INIT => "0000001000001110111000101000000010000010100001101010001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000001000000000001000000000000000000000000000000000000000000000000010000000100000000000000000000000") port map( O =>C_47_S_0_L_6_out, I0 =>  inp_feat(362), I1 =>  inp_feat(445), I2 =>  inp_feat(384), I3 =>  inp_feat(284), I4 =>  inp_feat(152), I5 =>  inp_feat(134), I6 =>  inp_feat(150), I7 =>  inp_feat(29)); 
C_47_S_0_L_7_inst : LUT8 generic map(INIT => "0000001000000000101100100010000000000000010000001111000101010000001000101001000000000000000000000000000000100000011100000000000000000000000000001000001100010000000000000000000001110100000000000000000000000000000000000000000000000100000000000000000000000000") port map( O =>C_47_S_0_L_7_out, I0 =>  inp_feat(420), I1 =>  inp_feat(464), I2 =>  inp_feat(253), I3 =>  inp_feat(171), I4 =>  inp_feat(452), I5 =>  inp_feat(273), I6 =>  inp_feat(446), I7 =>  inp_feat(487)); 
C_47_S_1_L_0_inst : LUT8 generic map(INIT => "0000000100010001000000000000000000000000000101010000000000000000000000010000000000000000000000000000000000000000000000000000000000000010110100110000000000000000100000001101110100000000000000000000000000000000000000000000000000000010000000000000000000000000") port map( O =>C_47_S_1_L_0_out, I0 =>  inp_feat(273), I1 =>  inp_feat(384), I2 =>  inp_feat(200), I3 =>  inp_feat(221), I4 =>  inp_feat(132), I5 =>  inp_feat(476), I6 =>  inp_feat(290), I7 =>  inp_feat(391)); 
C_47_S_1_L_1_inst : LUT8 generic map(INIT => "0000010100010001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111101000000000000000000010000000000010000000000000000000000010101000100010000000000000001000100000000000000000000000000000") port map( O =>C_47_S_1_L_1_out, I0 =>  inp_feat(419), I1 =>  inp_feat(20), I2 =>  inp_feat(448), I3 =>  inp_feat(383), I4 =>  inp_feat(68), I5 =>  inp_feat(487), I6 =>  inp_feat(242), I7 =>  inp_feat(235)); 
C_47_S_1_L_2_inst : LUT8 generic map(INIT => "1100101000100000000000000000001010001010100010010000000000100000101000001000000000000000100000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_47_S_1_L_2_out, I0 =>  inp_feat(217), I1 =>  inp_feat(207), I2 =>  inp_feat(475), I3 =>  inp_feat(265), I4 =>  inp_feat(102), I5 =>  inp_feat(494), I6 =>  inp_feat(31), I7 =>  inp_feat(172)); 
C_47_S_1_L_3_inst : LUT8 generic map(INIT => "1000001010110010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_1_L_3_out, I0 =>  inp_feat(172), I1 =>  inp_feat(142), I2 =>  inp_feat(32), I3 =>  inp_feat(81), I4 =>  inp_feat(93), I5 =>  inp_feat(251), I6 =>  inp_feat(49), I7 =>  inp_feat(242)); 
C_47_S_1_L_4_inst : LUT8 generic map(INIT => "0100000000000000010010000000000000000000000000000000010000000000111011000000000111011101000000000000000000000000010001011101010000000000000000000000000000000000000000000000000000000000000000000101000000000000110100000100010000000000000000000100000000000000") port map( O =>C_47_S_1_L_4_out, I0 =>  inp_feat(445), I1 =>  inp_feat(487), I2 =>  inp_feat(410), I3 =>  inp_feat(116), I4 =>  inp_feat(464), I5 =>  inp_feat(387), I6 =>  inp_feat(316), I7 =>  inp_feat(446)); 
C_47_S_1_L_5_inst : LUT8 generic map(INIT => "1111010101110100111111010000000100000000001000001000000000000000000000000000000010000000000000000000100000000000000000000000000001010101000000001000110101000111000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_1_L_5_out, I0 =>  inp_feat(73), I1 =>  inp_feat(291), I2 =>  inp_feat(244), I3 =>  inp_feat(373), I4 =>  inp_feat(204), I5 =>  inp_feat(296), I6 =>  inp_feat(446), I7 =>  inp_feat(37)); 
C_47_S_1_L_6_inst : LUT8 generic map(INIT => "1100100000001000000100000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_1_L_6_out, I0 =>  inp_feat(419), I1 =>  inp_feat(87), I2 =>  inp_feat(510), I3 =>  inp_feat(287), I4 =>  inp_feat(23), I5 =>  inp_feat(198), I6 =>  inp_feat(306), I7 =>  inp_feat(122)); 
C_47_S_1_L_7_inst : LUT8 generic map(INIT => "0100000100101001000000000000010100000000000000010000000000000001000111000100001000000000000000000000100010110011000000000000000011000100100010100000011100000100000010100000001100000000000000000000000000000001000000100000000100000000000000000000000000000001") port map( O =>C_47_S_1_L_7_out, I0 =>  inp_feat(445), I1 =>  inp_feat(229), I2 =>  inp_feat(301), I3 =>  inp_feat(504), I4 =>  inp_feat(294), I5 =>  inp_feat(207), I6 =>  inp_feat(457), I7 =>  inp_feat(304)); 
C_47_S_2_L_0_inst : LUT8 generic map(INIT => "0000010001001100000000000000000000000000010000000000000000000000000000001000000000001000100000000000000000000000000000000000000011011100110011000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_2_L_0_out, I0 =>  inp_feat(450), I1 =>  inp_feat(87), I2 =>  inp_feat(304), I3 =>  inp_feat(31), I4 =>  inp_feat(172), I5 =>  inp_feat(388), I6 =>  inp_feat(446), I7 =>  inp_feat(235)); 
C_47_S_2_L_1_inst : LUT8 generic map(INIT => "0011010101000000010111001000010000010000000000000000000000000000010000000000000010000000100000000101000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000") port map( O =>C_47_S_2_L_1_out, I0 =>  inp_feat(448), I1 =>  inp_feat(504), I2 =>  inp_feat(180), I3 =>  inp_feat(242), I4 =>  inp_feat(320), I5 =>  inp_feat(105), I6 =>  inp_feat(98), I7 =>  inp_feat(306)); 
C_47_S_2_L_2_inst : LUT8 generic map(INIT => "0000110001000000000000000000000000000000000000000000000000000000010011011001000000000001000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000110100000001000000000000000000001001000000000000000000000000") port map( O =>C_47_S_2_L_2_out, I0 =>  inp_feat(244), I1 =>  inp_feat(81), I2 =>  inp_feat(187), I3 =>  inp_feat(242), I4 =>  inp_feat(66), I5 =>  inp_feat(306), I6 =>  inp_feat(450), I7 =>  inp_feat(352)); 
C_47_S_2_L_3_inst : LUT8 generic map(INIT => "0110111100000000001110110000100000001001000010010000100000000000001110010000000000001000000010000000100000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_2_L_3_out, I0 =>  inp_feat(419), I1 =>  inp_feat(448), I2 =>  inp_feat(316), I3 =>  inp_feat(444), I4 =>  inp_feat(103), I5 =>  inp_feat(446), I6 =>  inp_feat(133), I7 =>  inp_feat(87)); 
C_47_S_2_L_4_inst : LUT8 generic map(INIT => "0000000010101000000000000000101000000000000000000000000000000000111000001010111000010000001000000000000010000000000000000000000000000000101010000000000000000000000000000000000000000000100010000000100010000000000000001000000000000000000000000000000000000000") port map( O =>C_47_S_2_L_4_out, I0 =>  inp_feat(469), I1 =>  inp_feat(411), I2 =>  inp_feat(494), I3 =>  inp_feat(221), I4 =>  inp_feat(81), I5 =>  inp_feat(114), I6 =>  inp_feat(273), I7 =>  inp_feat(20)); 
C_47_S_2_L_5_inst : LUT8 generic map(INIT => "0110100010001110000000000000100000000000000010000000000000001000000010000000100000100000000000000000000000000000000010000000000000001000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_2_L_5_out, I0 =>  inp_feat(229), I1 =>  inp_feat(485), I2 =>  inp_feat(20), I3 =>  inp_feat(464), I4 =>  inp_feat(287), I5 =>  inp_feat(116), I6 =>  inp_feat(126), I7 =>  inp_feat(81)); 
C_47_S_2_L_6_inst : LUT8 generic map(INIT => "0010001100000001001001110000010000000000000000000001010100000000000000000000000000110000000000100000000000000000000000000000000000000010000000001011001100010000000001000000000000001001000000000000000000000000000010000000000000000000000000000000000000000000") port map( O =>C_47_S_2_L_6_out, I0 =>  inp_feat(86), I1 =>  inp_feat(484), I2 =>  inp_feat(273), I3 =>  inp_feat(446), I4 =>  inp_feat(211), I5 =>  inp_feat(171), I6 =>  inp_feat(387), I7 =>  inp_feat(244)); 
C_47_S_2_L_7_inst : LUT8 generic map(INIT => "1101001100000000000000000000000010000000001000000010000000000000011011000000000010100000001000001000000000000000000000000000000011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_2_L_7_out, I0 =>  inp_feat(457), I1 =>  inp_feat(373), I2 =>  inp_feat(29), I3 =>  inp_feat(186), I4 =>  inp_feat(140), I5 =>  inp_feat(182), I6 =>  inp_feat(32), I7 =>  inp_feat(417)); 
C_47_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000010000000000100000110000001000100010110000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_3_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(51), I2 =>  inp_feat(478), I3 =>  inp_feat(378), I4 =>  inp_feat(207), I5 =>  inp_feat(36), I6 =>  inp_feat(132), I7 =>  inp_feat(87)); 
C_47_S_3_L_1_inst : LUT8 generic map(INIT => "1110001011010000100010100000000001000000111100000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_3_L_1_out, I0 =>  inp_feat(266), I1 =>  inp_feat(41), I2 =>  inp_feat(193), I3 =>  inp_feat(10), I4 =>  inp_feat(172), I5 =>  inp_feat(107), I6 =>  inp_feat(336), I7 =>  inp_feat(87)); 
C_47_S_3_L_2_inst : LUT8 generic map(INIT => "0001111100000111000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000001000010000000000000011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_3_L_2_out, I0 =>  inp_feat(204), I1 =>  inp_feat(473), I2 =>  inp_feat(179), I3 =>  inp_feat(325), I4 =>  inp_feat(290), I5 =>  inp_feat(407), I6 =>  inp_feat(132), I7 =>  inp_feat(380)); 
C_47_S_3_L_3_inst : LUT8 generic map(INIT => "1100000010110010011010000000000010000000100000000000000000000000100100001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_47_S_3_L_3_out, I0 =>  inp_feat(444), I1 =>  inp_feat(302), I2 =>  inp_feat(94), I3 =>  inp_feat(457), I4 =>  inp_feat(407), I5 =>  inp_feat(135), I6 =>  inp_feat(417), I7 =>  inp_feat(338)); 
C_47_S_3_L_4_inst : LUT8 generic map(INIT => "1010100000000000000000010000000000101010001000001001001100000010000010001000000000000000000000000000101100000000000000110000001100000000000000000000000000000000000000000000000000010001000000010000000000000000000000000000000000000000000000000000000000000010") port map( O =>C_47_S_3_L_4_out, I0 =>  inp_feat(388), I1 =>  inp_feat(372), I2 =>  inp_feat(50), I3 =>  inp_feat(446), I4 =>  inp_feat(274), I5 =>  inp_feat(445), I6 =>  inp_feat(442), I7 =>  inp_feat(116)); 
C_47_S_3_L_5_inst : LUT8 generic map(INIT => "0001000001010000000000000000000000100000001010000000000000000000000000000001000000000000000000001000100000100000000000000000000011010000001000000000000000000000110100001000101000101000101010100000000000110000000000000000000000000000101000100010000000100000") port map( O =>C_47_S_3_L_5_out, I0 =>  inp_feat(31), I1 =>  inp_feat(504), I2 =>  inp_feat(278), I3 =>  inp_feat(229), I4 =>  inp_feat(100), I5 =>  inp_feat(506), I6 =>  inp_feat(207), I7 =>  inp_feat(36)); 
C_47_S_3_L_6_inst : LUT8 generic map(INIT => "0101000111000001000000000000000000000000000000000000000000000000000011010100101100000000010000000000000000000000000000000000000001011010000000000000101000000000000000000000000000101010100000100000000001000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_3_L_6_out, I0 =>  inp_feat(134), I1 =>  inp_feat(179), I2 =>  inp_feat(364), I3 =>  inp_feat(475), I4 =>  inp_feat(444), I5 =>  inp_feat(172), I6 =>  inp_feat(86), I7 =>  inp_feat(272)); 
C_47_S_3_L_7_inst : LUT8 generic map(INIT => "0100010100000000000000000010000011000101010001000000011011000101101000000000000000000000001000000010000010000000011001000110010000000000000000000000000100000000110000000100110000000100100001000000000000000000000000000000000000000000000000000000000000000001") port map( O =>C_47_S_3_L_7_out, I0 =>  inp_feat(452), I1 =>  inp_feat(444), I2 =>  inp_feat(367), I3 =>  inp_feat(509), I4 =>  inp_feat(302), I5 =>  inp_feat(52), I6 =>  inp_feat(171), I7 =>  inp_feat(387)); 
C_47_S_4_L_0_inst : LUT8 generic map(INIT => "0100010100000000000000000000000000000000000000001100100000000000110111010000000010000100000000000000010000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_4_L_0_out, I0 =>  inp_feat(176), I1 =>  inp_feat(407), I2 =>  inp_feat(57), I3 =>  inp_feat(132), I4 =>  inp_feat(398), I5 =>  inp_feat(408), I6 =>  inp_feat(378), I7 =>  inp_feat(465)); 
C_47_S_4_L_1_inst : LUT8 generic map(INIT => "1111010100000001000000000000000000010000000100010000000100000000111100001001000000110000000000000001000010010000001000000000000000000001001000110000000000000000000000000010000000000000000000000000000000000000000100000001000100010000001000000010000000000000") port map( O =>C_47_S_4_L_1_out, I0 =>  inp_feat(204), I1 =>  inp_feat(61), I2 =>  inp_feat(407), I3 =>  inp_feat(264), I4 =>  inp_feat(455), I5 =>  inp_feat(207), I6 =>  inp_feat(457), I7 =>  inp_feat(465)); 
C_47_S_4_L_2_inst : LUT8 generic map(INIT => "0000010101000100010001000100000010000100000000000000000001000100000001000100010000000100000000000000000000000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_4_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(87), I2 =>  inp_feat(298), I3 =>  inp_feat(133), I4 =>  inp_feat(5), I5 =>  inp_feat(410), I6 =>  inp_feat(442), I7 =>  inp_feat(353)); 
C_47_S_4_L_3_inst : LUT8 generic map(INIT => "0000010000000000000000000000000010001000000000000000000000000000100110000000000000001000000000000000000000000000000000000000000011000110001001000010000000000000100000100111010000000010000000001100000001000000000000000000000001000000000000000000000000000000") port map( O =>C_47_S_4_L_3_out, I0 =>  inp_feat(302), I1 =>  inp_feat(413), I2 =>  inp_feat(457), I3 =>  inp_feat(278), I4 =>  inp_feat(217), I5 =>  inp_feat(475), I6 =>  inp_feat(31), I7 =>  inp_feat(247)); 
C_47_S_4_L_4_inst : LUT8 generic map(INIT => "1000000000000000101010000000000000101110000000100000000000000000000000000000000000000000000000000010000000000000000000000000000011100000100000001010000010100000101000000010000010100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_4_L_4_out, I0 =>  inp_feat(407), I1 =>  inp_feat(134), I2 =>  inp_feat(336), I3 =>  inp_feat(278), I4 =>  inp_feat(384), I5 =>  inp_feat(406), I6 =>  inp_feat(34), I7 =>  inp_feat(316)); 
C_47_S_4_L_5_inst : LUT8 generic map(INIT => "0001110011110100100100001011000000110000001100000000000000110000000000000010000000100000001000000011000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_47_S_4_L_5_out, I0 =>  inp_feat(445), I1 =>  inp_feat(316), I2 =>  inp_feat(336), I3 =>  inp_feat(179), I4 =>  inp_feat(31), I5 =>  inp_feat(490), I6 =>  inp_feat(444), I7 =>  inp_feat(438)); 
C_47_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000101000000010000010100000000000001010000000000000001000000001000010000000000000001010001001000000101000000000000010100000000000101011000000000000000000000000000000000000000000000010000010000010100000000100001000000000000000000000000000000000") port map( O =>C_47_S_4_L_6_out, I0 =>  inp_feat(217), I1 =>  inp_feat(61), I2 =>  inp_feat(455), I3 =>  inp_feat(207), I4 =>  inp_feat(73), I5 =>  inp_feat(384), I6 =>  inp_feat(457), I7 =>  inp_feat(171)); 
C_47_S_4_L_7_inst : LUT8 generic map(INIT => "0010101000101010011000110010100000000010000000000000000000001011001000100000101000000010000010100000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000001000000000000000100000000000000000000010000000001000000000") port map( O =>C_47_S_4_L_7_out, I0 =>  inp_feat(287), I1 =>  inp_feat(452), I2 =>  inp_feat(134), I3 =>  inp_feat(410), I4 =>  inp_feat(402), I5 =>  inp_feat(486), I6 =>  inp_feat(133), I7 =>  inp_feat(446)); 
C_48_S_0_L_0_inst : LUT8 generic map(INIT => "1111111111111111111110110000000011011010010100011000101000000000100010001001000010001000000000000100000000000000000000000000000010100010111111000010001000000000100000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_48_S_0_L_0_out, I0 =>  inp_feat(153), I1 =>  inp_feat(272), I2 =>  inp_feat(373), I3 =>  inp_feat(155), I4 =>  inp_feat(229), I5 =>  inp_feat(54), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_48_S_0_L_1_inst : LUT8 generic map(INIT => "1110110011001100101010000000111111001100110011000000100000000000101011111000100000000000000010111111111110001000000000000000000011001110110011001100111100001010100010000100110000000000000000001000101000001000001010100000100000001100000010000000100000000000") port map( O =>C_48_S_0_L_1_out, I0 =>  inp_feat(267), I1 =>  inp_feat(87), I2 =>  inp_feat(340), I3 =>  inp_feat(46), I4 =>  inp_feat(310), I5 =>  inp_feat(56), I6 =>  inp_feat(256), I7 =>  inp_feat(71)); 
C_48_S_0_L_2_inst : LUT8 generic map(INIT => "1010100011111000101110101000101010111000011100001010100010000000110010000000100010000000000000001001000000000000011100000000000011111110111010101001000010101000111110001010101000000000000000000000100000001000000000000000000010010000000000000001000000000000") port map( O =>C_48_S_0_L_2_out, I0 =>  inp_feat(224), I1 =>  inp_feat(370), I2 =>  inp_feat(54), I3 =>  inp_feat(139), I4 =>  inp_feat(183), I5 =>  inp_feat(71), I6 =>  inp_feat(151), I7 =>  inp_feat(266)); 
C_48_S_0_L_3_inst : LUT8 generic map(INIT => "1110110110000000110000000000000011111011101100100000000000000000011110001000100001000000000000001011000110101010000000100010100011111000101010001111000010100000101010001010000000000000001000000000000000000000000000001010000000100000001000000000000010000000") port map( O =>C_48_S_0_L_3_out, I0 =>  inp_feat(427), I1 =>  inp_feat(166), I2 =>  inp_feat(504), I3 =>  inp_feat(266), I4 =>  inp_feat(296), I5 =>  inp_feat(135), I6 =>  inp_feat(183), I7 =>  inp_feat(311)); 
C_48_S_0_L_4_inst : LUT8 generic map(INIT => "0001101011101010100010001000101011101110100010101000100010001010110110101000101000000000110011101110111001111111000000110000111011100000101000101100000000000010101000000000100000000000000000001110000000000000010000000000000000100010000000000000000000000000") port map( O =>C_48_S_0_L_4_out, I0 =>  inp_feat(384), I1 =>  inp_feat(373), I2 =>  inp_feat(435), I3 =>  inp_feat(396), I4 =>  inp_feat(439), I5 =>  inp_feat(475), I6 =>  inp_feat(183), I7 =>  inp_feat(311)); 
C_48_S_0_L_5_inst : LUT8 generic map(INIT => "1111011011000000111100001010000011111000011000101111000011110010111111111011000011110000111000001111100000101000111100001110101001100100010000000010000010000000111010000000000011100000110000001111000110100000111100001110000011111000101000001110000010110000") port map( O =>C_48_S_0_L_5_out, I0 =>  inp_feat(120), I1 =>  inp_feat(373), I2 =>  inp_feat(267), I3 =>  inp_feat(105), I4 =>  inp_feat(282), I5 =>  inp_feat(221), I6 =>  inp_feat(340), I7 =>  inp_feat(74)); 
C_48_S_0_L_6_inst : LUT8 generic map(INIT => "1111111000001100111011001000110011010100010001001000010001001100111000000000010011000000100000001110000000000000011100000000000010101010000010001000110000000000000000000000000000000000000000001010001000000000101000001000000000000000000000000000000000000000") port map( O =>C_48_S_0_L_6_out, I0 =>  inp_feat(6), I1 =>  inp_feat(183), I2 =>  inp_feat(191), I3 =>  inp_feat(60), I4 =>  inp_feat(416), I5 =>  inp_feat(483), I6 =>  inp_feat(92), I7 =>  inp_feat(296)); 
C_48_S_0_L_7_inst : LUT8 generic map(INIT => "1100101000001010011110101000101000001010000010101100101010001010111010100000100011001000001010001010000000000000100000000000100011000000000000001100000010000000110000000010001010001000000010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_48_S_0_L_7_out, I0 =>  inp_feat(459), I1 =>  inp_feat(342), I2 =>  inp_feat(46), I3 =>  inp_feat(291), I4 =>  inp_feat(364), I5 =>  inp_feat(266), I6 =>  inp_feat(285), I7 =>  inp_feat(33)); 
C_48_S_1_L_0_inst : LUT8 generic map(INIT => "1111111111100010001111110010000011110000111100100101001000110000111011101010101011101010001000001111101001100010111100000000000011010101100000000101001000000000111100111100010001010000000000001011000010000000011100000000000011100000110000000011000000000000") port map( O =>C_48_S_1_L_0_out, I0 =>  inp_feat(467), I1 =>  inp_feat(298), I2 =>  inp_feat(183), I3 =>  inp_feat(259), I4 =>  inp_feat(87), I5 =>  inp_feat(340), I6 =>  inp_feat(115), I7 =>  inp_feat(160)); 
C_48_S_1_L_1_inst : LUT8 generic map(INIT => "1110100011101010001010001100000011101000100010101100000011000000101010101000100010110010101000100000100000000000000000000000000000101000111010001000100011001010110011000000000011001100110011001010101010100010101010001010001010101000101000001010001010100000") port map( O =>C_48_S_1_L_1_out, I0 =>  inp_feat(54), I1 =>  inp_feat(87), I2 =>  inp_feat(428), I3 =>  inp_feat(317), I4 =>  inp_feat(387), I5 =>  inp_feat(130), I6 =>  inp_feat(492), I7 =>  inp_feat(11)); 
C_48_S_1_L_2_inst : LUT8 generic map(INIT => "1111111011101110101100000011000011110000100010111011000000000000111011001000101001100000001000001100000010000000000000000000000010101010101010101010000010100010100000000000000000000000000000001010001010001010100000000000000000000000000000000000000000000000") port map( O =>C_48_S_1_L_2_out, I0 =>  inp_feat(439), I1 =>  inp_feat(373), I2 =>  inp_feat(210), I3 =>  inp_feat(71), I4 =>  inp_feat(306), I5 =>  inp_feat(398), I6 =>  inp_feat(316), I7 =>  inp_feat(95)); 
C_48_S_1_L_3_inst : LUT8 generic map(INIT => "1110111011111000111110101110010001100000111010001111100011001000100010001110101011100000110010001000000011101010010000000100000001001101000010001111100011101000000000000000000000000000000000001010100010101010101010101010100000000000010000000000000000000000") port map( O =>C_48_S_1_L_3_out, I0 =>  inp_feat(387), I1 =>  inp_feat(87), I2 =>  inp_feat(183), I3 =>  inp_feat(277), I4 =>  inp_feat(340), I5 =>  inp_feat(259), I6 =>  inp_feat(412), I7 =>  inp_feat(216)); 
C_48_S_1_L_4_inst : LUT8 generic map(INIT => "1000101011101010001000001000000000101000110011101010100000001000110011000000100000001000000000001100100000001000000010000000000010000010100010101010100010000000000010100000101000001010000010101000101000000010000010000000000000001010000010000000100000001010") port map( O =>C_48_S_1_L_4_out, I0 =>  inp_feat(466), I1 =>  inp_feat(310), I2 =>  inp_feat(169), I3 =>  inp_feat(316), I4 =>  inp_feat(149), I5 =>  inp_feat(221), I6 =>  inp_feat(95), I7 =>  inp_feat(385)); 
C_48_S_1_L_5_inst : LUT8 generic map(INIT => "0110101001000111000111110000001011101111110111110111111100000100000010000000100001011111000000001100100001001100111111010000010011111111101011110011001100010001000001010101110101110101010101010101111101011111001100110100000001000000010101010101010100000101") port map( O =>C_48_S_1_L_5_out, I0 =>  inp_feat(56), I1 =>  inp_feat(263), I2 =>  inp_feat(64), I3 =>  inp_feat(33), I4 =>  inp_feat(285), I5 =>  inp_feat(282), I6 =>  inp_feat(90), I7 =>  inp_feat(266)); 
C_48_S_1_L_6_inst : LUT8 generic map(INIT => "1111010011000100111110001100110011101000000000000000100000000000011000000000000000000000101000001100000000000000000000000000000011010110110001011111111110000000000010000000000000000000000000000010100010101000000000000000000000000000000000000000000000000000") port map( O =>C_48_S_1_L_6_out, I0 =>  inp_feat(238), I1 =>  inp_feat(183), I2 =>  inp_feat(365), I3 =>  inp_feat(80), I4 =>  inp_feat(179), I5 =>  inp_feat(191), I6 =>  inp_feat(349), I7 =>  inp_feat(449)); 
C_48_S_1_L_7_inst : LUT8 generic map(INIT => "0100010111011101110011100000110001011101111111101100110010000100110011001110110011001100110011001100111011111100100011001000110001011010000000000000101000000000000011010000000000000000000000000000100000000000000000100000000001000100000000000000000000000000") port map( O =>C_48_S_1_L_7_out, I0 =>  inp_feat(328), I1 =>  inp_feat(428), I2 =>  inp_feat(221), I3 =>  inp_feat(142), I4 =>  inp_feat(42), I5 =>  inp_feat(316), I6 =>  inp_feat(500), I7 =>  inp_feat(266)); 
C_48_S_2_L_0_inst : LUT8 generic map(INIT => "1110101011101010111000101110001011101010111010101100010011000010100000001110100001111011110111111110100011101010110011001110111100000000110000001010111001001010111000000100000001000101000001001100110000000001111011110100111111000000000011000100110101001111") port map( O =>C_48_S_2_L_0_out, I0 =>  inp_feat(285), I1 =>  inp_feat(268), I2 =>  inp_feat(282), I3 =>  inp_feat(473), I4 =>  inp_feat(302), I5 =>  inp_feat(378), I6 =>  inp_feat(200), I7 =>  inp_feat(71)); 
C_48_S_2_L_1_inst : LUT8 generic map(INIT => "1110100011111111010111100101110110000000001010100000100000000000100010001111110111111000111101011000100010001100100010000000000001100010010010101111000001100110000000101000101000001000000000000000000011011101010000000101010100000000000010000000000000000000") port map( O =>C_48_S_2_L_1_out, I0 =>  inp_feat(15), I1 =>  inp_feat(451), I2 =>  inp_feat(327), I3 =>  inp_feat(221), I4 =>  inp_feat(212), I5 =>  inp_feat(385), I6 =>  inp_feat(378), I7 =>  inp_feat(71)); 
C_48_S_2_L_2_inst : LUT8 generic map(INIT => "1110110010100000101000001010000011111111000000001010111111110111111110001000100010000000100000000011000000000000101000100000001011001011000000001010000010100000001010000000000010100010101000101100100010000000101010001010000000100000000000001010001011101010") port map( O =>C_48_S_2_L_2_out, I0 =>  inp_feat(87), I1 =>  inp_feat(428), I2 =>  inp_feat(365), I3 =>  inp_feat(1), I4 =>  inp_feat(194), I5 =>  inp_feat(370), I6 =>  inp_feat(103), I7 =>  inp_feat(12)); 
C_48_S_2_L_3_inst : LUT8 generic map(INIT => "0110100010101010111100111100101010100000101000001100000000000000111000001000101011100000001000001000000000000000000000000000000010010010000000001100101010000010000000000000000011000010000000001110101000100000111000100000000000100010000000000000000000000000") port map( O =>C_48_S_2_L_3_out, I0 =>  inp_feat(206), I1 =>  inp_feat(41), I2 =>  inp_feat(310), I3 =>  inp_feat(285), I4 =>  inp_feat(100), I5 =>  inp_feat(267), I6 =>  inp_feat(151), I7 =>  inp_feat(437)); 
C_48_S_2_L_4_inst : LUT8 generic map(INIT => "1111110011100110111011110000011011001100101011101111101010000011111011100010001010101111000010100000000000000010101111110000001011001100000000000111001000001100110111100000000000000000010000001111111001110111111111110011011100000000000000000000101000000000") port map( O =>C_48_S_2_L_4_out, I0 =>  inp_feat(365), I1 =>  inp_feat(103), I2 =>  inp_feat(15), I3 =>  inp_feat(201), I4 =>  inp_feat(329), I5 =>  inp_feat(90), I6 =>  inp_feat(130), I7 =>  inp_feat(323)); 
C_48_S_2_L_5_inst : LUT8 generic map(INIT => "1110110010001101110011001100010011000100000000000000010000000000111111001000111110001000100011011111111100000000000000010000000111101100000001000100010000001000010001000000000000000100000000000000000000000000000000000000110000000000000000000000000000000001") port map( O =>C_48_S_2_L_5_out, I0 =>  inp_feat(265), I1 =>  inp_feat(296), I2 =>  inp_feat(107), I3 =>  inp_feat(224), I4 =>  inp_feat(370), I5 =>  inp_feat(495), I6 =>  inp_feat(311), I7 =>  inp_feat(183)); 
C_48_S_2_L_6_inst : LUT8 generic map(INIT => "1101100011001000001000001111000011001000110010001111000011110000111101000010000001000000100000001000100000000000110000001000000001110101111100001000000010000000001000001010100011110000111000001101000000000000000000000000000000001000000000000110000010000000") port map( O =>C_48_S_2_L_6_out, I0 =>  inp_feat(214), I1 =>  inp_feat(33), I2 =>  inp_feat(229), I3 =>  inp_feat(65), I4 =>  inp_feat(381), I5 =>  inp_feat(302), I6 =>  inp_feat(218), I7 =>  inp_feat(272)); 
C_48_S_2_L_7_inst : LUT8 generic map(INIT => "1111011111111110101100101010000011110010111000100100000011110010101101101111111100100000000000001111000011001000101000001101000011111011111111101010000011110000101000101011101011110011111100101111101011111010001000001111000111110010111110001010000011110100") port map( O =>C_48_S_2_L_7_out, I0 =>  inp_feat(103), I1 =>  inp_feat(317), I2 =>  inp_feat(87), I3 =>  inp_feat(101), I4 =>  inp_feat(33), I5 =>  inp_feat(56), I6 =>  inp_feat(203), I7 =>  inp_feat(64)); 
C_48_S_3_L_0_inst : LUT8 generic map(INIT => "1111100011010101111100001111000000001000110101001100000011000000100010000000000011011101111110000000000000000000000010000000000010110000101000001011000011000000000000000000000000000000000000001111100010100010000000101111101000000000000000000000000000000000") port map( O =>C_48_S_3_L_0_out, I0 =>  inp_feat(365), I1 =>  inp_feat(229), I2 =>  inp_feat(267), I3 =>  inp_feat(422), I4 =>  inp_feat(288), I5 =>  inp_feat(466), I6 =>  inp_feat(109), I7 =>  inp_feat(437)); 
C_48_S_3_L_1_inst : LUT8 generic map(INIT => "0011010011101100111101101110000010100001000110000100000100010000111110011111101010110011101000100110111101010000001100100000000011010000010000001101110001000000110000000000000011000100000000001100000011000000000000000000000000000000000000001000000000000000") port map( O =>C_48_S_3_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(383), I2 =>  inp_feat(310), I3 =>  inp_feat(210), I4 =>  inp_feat(340), I5 =>  inp_feat(267), I6 =>  inp_feat(151), I7 =>  inp_feat(378)); 
C_48_S_3_L_2_inst : LUT8 generic map(INIT => "1111111011111111101010001011111110111000101110100010111000111111111111001101110001110100001111010110010011110100011011110010110101011110110001101110111010101101100101000000000000000000001011111010100001000100100011110001110101000101000000000100010100001100") port map( O =>C_48_S_3_L_2_out, I0 =>  inp_feat(329), I1 =>  inp_feat(108), I2 =>  inp_feat(282), I3 =>  inp_feat(473), I4 =>  inp_feat(101), I5 =>  inp_feat(130), I6 =>  inp_feat(218), I7 =>  inp_feat(272)); 
C_48_S_3_L_3_inst : LUT8 generic map(INIT => "1111111100010101110111111111000011001111101000001100111000000000110011110101111111001111100000000000010000000000000001000000000011101001100010111100111100000001110011110000001011001110000000100000000110000010010000010001000100000000000000000000000000000000") port map( O =>C_48_S_3_L_3_out, I0 =>  inp_feat(107), I1 =>  inp_feat(307), I2 =>  inp_feat(338), I3 =>  inp_feat(504), I4 =>  inp_feat(340), I5 =>  inp_feat(238), I6 =>  inp_feat(267), I7 =>  inp_feat(151)); 
C_48_S_3_L_4_inst : LUT8 generic map(INIT => "1001010011100110111001110000010001101110110001100010010011001100111101101010000010110000000000000000000000100010001000100000000010101110101000100010001000000000001000101010001000100010000000001010000000000000001000000000000000000000000000000010000000000000") port map( O =>C_48_S_3_L_4_out, I0 =>  inp_feat(380), I1 =>  inp_feat(128), I2 =>  inp_feat(298), I3 =>  inp_feat(214), I4 =>  inp_feat(468), I5 =>  inp_feat(267), I6 =>  inp_feat(210), I7 =>  inp_feat(151)); 
C_48_S_3_L_5_inst : LUT8 generic map(INIT => "1100110101101100111110111000110011011111101011101100110010101110011111011010111001010000001011101110110000001110010000001010101010111011101010101010000000100010000111010000110000000100000001000011011100001000001000000000101000111101101011100000010000100000") port map( O =>C_48_S_3_L_5_out, I0 =>  inp_feat(15), I1 =>  inp_feat(382), I2 =>  inp_feat(221), I3 =>  inp_feat(56), I4 =>  inp_feat(331), I5 =>  inp_feat(328), I6 =>  inp_feat(71), I7 =>  inp_feat(152)); 
C_48_S_3_L_6_inst : LUT8 generic map(INIT => "1111111111111111111000011010101010110010101110101000000010101010111100011011000010000000000000101001000010110000100000000000000001111110111111111110001110001000100000001011100010000000100010100001100000110000000000000000000000100000101100001000000010001000") port map( O =>C_48_S_3_L_6_out, I0 =>  inp_feat(42), I1 =>  inp_feat(105), I2 =>  inp_feat(373), I3 =>  inp_feat(340), I4 =>  inp_feat(310), I5 =>  inp_feat(370), I6 =>  inp_feat(507), I7 =>  inp_feat(71)); 
C_48_S_3_L_7_inst : LUT8 generic map(INIT => "1111100011110000101100001011100011111110111100000101010000000000111111111010001011110111100000001111011000101010000000100000000011010010100100000001000000001000100000000000000000000000000000000101101000000000000000000000000011111000000000000000000000000000") port map( O =>C_48_S_3_L_7_out, I0 =>  inp_feat(428), I1 =>  inp_feat(149), I2 =>  inp_feat(54), I3 =>  inp_feat(183), I4 =>  inp_feat(87), I5 =>  inp_feat(33), I6 =>  inp_feat(1), I7 =>  inp_feat(58)); 
C_48_S_4_L_0_inst : LUT8 generic map(INIT => "0110010010101000111010101010000011101110101010101010101010111001101010001010100010101000100010001000101000100000100000001010000011111101101110001011100010110010111111111010101101010000110100001010000000100000000000000011000010101010001100000010000000010000") port map( O =>C_48_S_4_L_0_out, I0 =>  inp_feat(267), I1 =>  inp_feat(296), I2 =>  inp_feat(58), I3 =>  inp_feat(509), I4 =>  inp_feat(183), I5 =>  inp_feat(31), I6 =>  inp_feat(238), I7 =>  inp_feat(262)); 
C_48_S_4_L_1_inst : LUT8 generic map(INIT => "1100111010101000111111011000111011101100100000001110010000000000111011001010111011111111101011101110000010100100000000000000000010100000001000000101000010110010000000001010000010100000101100001010000000000000101100101010001010100000101000001010000010110000") port map( O =>C_48_S_4_L_1_out, I0 =>  inp_feat(365), I1 =>  inp_feat(268), I2 =>  inp_feat(87), I3 =>  inp_feat(101), I4 =>  inp_feat(329), I5 =>  inp_feat(130), I6 =>  inp_feat(64), I7 =>  inp_feat(33)); 
C_48_S_4_L_2_inst : LUT8 generic map(INIT => "1111111111001010100011100010101011001110000011100000110110001001010001111100111100000000000000100000100000001010000000000000000011001110100011001010111110101010110011101000101011001111100010111100111011111010000010110000001000000000000010110000000000000000") port map( O =>C_48_S_4_L_2_out, I0 =>  inp_feat(108), I1 =>  inp_feat(54), I2 =>  inp_feat(200), I3 =>  inp_feat(90), I4 =>  inp_feat(392), I5 =>  inp_feat(33), I6 =>  inp_feat(87), I7 =>  inp_feat(64)); 
C_48_S_4_L_3_inst : LUT8 generic map(INIT => "1100100011111000010010000111000000000000111100000000000001010000111110000000000011001000000000001100000000000000000000000000000011001000110011001000000010000000110000000100000000000000100000000000000000000000100000001000000011000000000000001100000010000000") port map( O =>C_48_S_4_L_3_out, I0 =>  inp_feat(200), I1 =>  inp_feat(392), I2 =>  inp_feat(486), I3 =>  inp_feat(444), I4 =>  inp_feat(297), I5 =>  inp_feat(428), I6 =>  inp_feat(288), I7 =>  inp_feat(435)); 
C_48_S_4_L_4_inst : LUT8 generic map(INIT => "0101001111111100110101000010000010000111011011100000000000000000110110011101010010001000000100000001010101000101000000000001000110111110000000000000111000000000101111100001000000000100000000000001110000000000000011000000000000010000000100000101110100010000") port map( O =>C_48_S_4_L_4_out, I0 =>  inp_feat(317), I1 =>  inp_feat(272), I2 =>  inp_feat(365), I3 =>  inp_feat(266), I4 =>  inp_feat(373), I5 =>  inp_feat(428), I6 =>  inp_feat(288), I7 =>  inp_feat(435)); 
C_48_S_4_L_5_inst : LUT8 generic map(INIT => "1000011001011101110010000010001011110010100110101000000000000000111011000111110010100010000000001010001010100000111000000000000010001111111111100010001000101010001110111001001000000000000000001111111111111110000000000000000001110100001100000000000000000000") port map( O =>C_48_S_4_L_5_out, I0 =>  inp_feat(297), I1 =>  inp_feat(176), I2 =>  inp_feat(210), I3 =>  inp_feat(412), I4 =>  inp_feat(282), I5 =>  inp_feat(255), I6 =>  inp_feat(340), I7 =>  inp_feat(433)); 
C_48_S_4_L_6_inst : LUT8 generic map(INIT => "1110100011001100110000000000000000101110010011001101010011111101110111001110010101000100111101001100110011010101110010001110010100000100000000000000000000000000010000000000000001010100111100001100110010100000110000001000000000000100000000001101010001110000") port map( O =>C_48_S_4_L_6_out, I0 =>  inp_feat(336), I1 =>  inp_feat(306), I2 =>  inp_feat(367), I3 =>  inp_feat(328), I4 =>  inp_feat(414), I5 =>  inp_feat(420), I6 =>  inp_feat(221), I7 =>  inp_feat(480)); 
C_48_S_4_L_7_inst : LUT8 generic map(INIT => "1010110011101110001000000010000000001000000010100000000000000000111111101010001000001100000000000000000000000010000000000000000010001000000000001010000010100000000010000000000000000000000000001010101000101010100010100010100000100010000010101000100000000000") port map( O =>C_48_S_4_L_7_out, I0 =>  inp_feat(296), I1 =>  inp_feat(53), I2 =>  inp_feat(221), I3 =>  inp_feat(316), I4 =>  inp_feat(42), I5 =>  inp_feat(1), I6 =>  inp_feat(81), I7 =>  inp_feat(282)); 
C_49_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000100000000000000000000000000000000010000000001000001000010000101110001011000100111000000000001000001010000001100000000000000000000000000000000001100000000000000010100001000000000000000100001001100000000001100010000000000000000000000000000000001") port map( O =>C_49_S_0_L_0_out, I0 =>  inp_feat(33), I1 =>  inp_feat(282), I2 =>  inp_feat(183), I3 =>  inp_feat(267), I4 =>  inp_feat(11), I5 =>  inp_feat(106), I6 =>  inp_feat(54), I7 =>  inp_feat(111)); 
C_49_S_0_L_1_inst : LUT8 generic map(INIT => "0010000000000010000000000000000010000011101000100100000011110101000000000000000000000000000000000000000000010000000000000001000000010000101110000001000011010001011100111010000001010111101100000000000000000000000000000001001000000000001000000001001000100000") port map( O =>C_49_S_0_L_1_out, I0 =>  inp_feat(154), I1 =>  inp_feat(11), I2 =>  inp_feat(340), I3 =>  inp_feat(267), I4 =>  inp_feat(216), I5 =>  inp_feat(71), I6 =>  inp_feat(266), I7 =>  inp_feat(160)); 
C_49_S_0_L_2_inst : LUT8 generic map(INIT => "1010000010100000100000001011101011110000001010100111000001110010000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000100000100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_0_L_2_out, I0 =>  inp_feat(328), I1 =>  inp_feat(380), I2 =>  inp_feat(409), I3 =>  inp_feat(221), I4 =>  inp_feat(331), I5 =>  inp_feat(390), I6 =>  inp_feat(305), I7 =>  inp_feat(294)); 
C_49_S_0_L_3_inst : LUT8 generic map(INIT => "0010101000100110101010100000101000100111000000011010101000000000000000100000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_0_L_3_out, I0 =>  inp_feat(210), I1 =>  inp_feat(413), I2 =>  inp_feat(373), I3 =>  inp_feat(328), I4 =>  inp_feat(213), I5 =>  inp_feat(111), I6 =>  inp_feat(322), I7 =>  inp_feat(305)); 
C_49_S_0_L_4_inst : LUT8 generic map(INIT => "1000000010001000001000000000001000000000000000000100000000100000101100001000000011101010001010001110000010000000010100000011100000000000000000000000100000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000") port map( O =>C_49_S_0_L_4_out, I0 =>  inp_feat(301), I1 =>  inp_feat(228), I2 =>  inp_feat(164), I3 =>  inp_feat(385), I4 =>  inp_feat(200), I5 =>  inp_feat(221), I6 =>  inp_feat(71), I7 =>  inp_feat(163)); 
C_49_S_0_L_5_inst : LUT8 generic map(INIT => "0111000000010001000001000000000000000000000000000111011100000000000101110111011100010111000000100000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000") port map( O =>C_49_S_0_L_5_out, I0 =>  inp_feat(216), I1 =>  inp_feat(387), I2 =>  inp_feat(428), I3 =>  inp_feat(291), I4 =>  inp_feat(15), I5 =>  inp_feat(106), I6 =>  inp_feat(108), I7 =>  inp_feat(322)); 
C_49_S_0_L_6_inst : LUT8 generic map(INIT => "0111000000010001001000001111000000010000001101110001000011111111000000000000000010101010100000000000000000111010100000001010101000000000000000000000000001000000000000000001010100000000011111000000000000000000000000000000000000000000000100010000000010111000") port map( O =>C_49_S_0_L_6_out, I0 =>  inp_feat(87), I1 =>  inp_feat(323), I2 =>  inp_feat(340), I3 =>  inp_feat(54), I4 =>  inp_feat(90), I5 =>  inp_feat(1), I6 =>  inp_feat(106), I7 =>  inp_feat(64)); 
C_49_S_0_L_7_inst : LUT8 generic map(INIT => "0000110011000100010101000111110001001100000000000001000100000001010001000000010100000101111001000000001000001011000001110000000100000000000000000000000001100000000000000000000000000000001000010000000000000000000000000000000000000011000100100000000000000000") port map( O =>C_49_S_0_L_7_out, I0 =>  inp_feat(71), I1 =>  inp_feat(362), I2 =>  inp_feat(483), I3 =>  inp_feat(331), I4 =>  inp_feat(1), I5 =>  inp_feat(329), I6 =>  inp_feat(390), I7 =>  inp_feat(163)); 
C_49_S_1_L_0_inst : LUT8 generic map(INIT => "0100000001000000010000001100000000000000000000000000000000000000000000001110010001000000010000000000000010000000100000001000000011000000010000000000000001000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000") port map( O =>C_49_S_1_L_0_out, I0 =>  inp_feat(310), I1 =>  inp_feat(435), I2 =>  inp_feat(151), I3 =>  inp_feat(183), I4 =>  inp_feat(60), I5 =>  inp_feat(266), I6 =>  inp_feat(102), I7 =>  inp_feat(160)); 
C_49_S_1_L_1_inst : LUT8 generic map(INIT => "0100110010110100000000000000000001000100110000001000000000000000000000001000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_1_L_1_out, I0 =>  inp_feat(385), I1 =>  inp_feat(219), I2 =>  inp_feat(459), I3 =>  inp_feat(471), I4 =>  inp_feat(409), I5 =>  inp_feat(1), I6 =>  inp_feat(500), I7 =>  inp_feat(305)); 
C_49_S_1_L_2_inst : LUT8 generic map(INIT => "1011001011110010010100000011001100000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_1_L_2_out, I0 =>  inp_feat(161), I1 =>  inp_feat(232), I2 =>  inp_feat(107), I3 =>  inp_feat(428), I4 =>  inp_feat(340), I5 =>  inp_feat(311), I6 =>  inp_feat(444), I7 =>  inp_feat(305)); 
C_49_S_1_L_3_inst : LUT8 generic map(INIT => "0011000010000010110111000000000000000000000100000101000000010000110100001010101011010000000000000000000010000000100100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_1_L_3_out, I0 =>  inp_feat(439), I1 =>  inp_feat(221), I2 =>  inp_feat(328), I3 =>  inp_feat(329), I4 =>  inp_feat(428), I5 =>  inp_feat(52), I6 =>  inp_feat(316), I7 =>  inp_feat(305)); 
C_49_S_1_L_4_inst : LUT8 generic map(INIT => "0011000000011000000000000000001001000000011101010100000000010000010000000000000000000000000000000000000000000000000000000000000011110111010100000011000000000011100100001101000000110000000000010000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_1_L_4_out, I0 =>  inp_feat(267), I1 =>  inp_feat(307), I2 =>  inp_feat(317), I3 =>  inp_feat(183), I4 =>  inp_feat(0), I5 =>  inp_feat(373), I6 =>  inp_feat(305), I7 =>  inp_feat(11)); 
C_49_S_1_L_5_inst : LUT8 generic map(INIT => "0010000000000000000000000000000010100000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000011111111001100000101000000000000101100000000000000000000000000001111111111011111000100000100000100000000000000000000000000000000") port map( O =>C_49_S_1_L_5_out, I0 =>  inp_feat(103), I1 =>  inp_feat(90), I2 =>  inp_feat(340), I3 =>  inp_feat(64), I4 =>  inp_feat(12), I5 =>  inp_feat(60), I6 =>  inp_feat(106), I7 =>  inp_feat(216)); 
C_49_S_1_L_6_inst : LUT8 generic map(INIT => "0111111000101110001000101000101100001000100010001000000000001000001011001000100000000000100010100000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000010100000010000000010000000100000000000000000000000000000000000000") port map( O =>C_49_S_1_L_6_out, I0 =>  inp_feat(383), I1 =>  inp_feat(198), I2 =>  inp_feat(373), I3 =>  inp_feat(183), I4 =>  inp_feat(216), I5 =>  inp_feat(214), I6 =>  inp_feat(259), I7 =>  inp_feat(288)); 
C_49_S_1_L_7_inst : LUT8 generic map(INIT => "0010000000000000000000000000000000000000000000000000000000000000101110001000000000000000000000001000000000000000010000000000000000000111100011000000001000000000000000000000000000000000000000000001110100000000000011010000000001000001000000000000000000000000") port map( O =>C_49_S_1_L_7_out, I0 =>  inp_feat(405), I1 =>  inp_feat(316), I2 =>  inp_feat(380), I3 =>  inp_feat(15), I4 =>  inp_feat(349), I5 =>  inp_feat(294), I6 =>  inp_feat(306), I7 =>  inp_feat(106)); 
C_49_S_2_L_0_inst : LUT8 generic map(INIT => "0000100001100000111010001100000000000000000000000100000000000000100000000100000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_2_L_0_out, I0 =>  inp_feat(154), I1 =>  inp_feat(143), I2 =>  inp_feat(239), I3 =>  inp_feat(266), I4 =>  inp_feat(267), I5 =>  inp_feat(12), I6 =>  inp_feat(89), I7 =>  inp_feat(305)); 
C_49_S_2_L_1_inst : LUT8 generic map(INIT => "1000000010000000000000000000000010100000101101001000000000000000000000001010000000000000100000001010000010111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_2_L_1_out, I0 =>  inp_feat(15), I1 =>  inp_feat(26), I2 =>  inp_feat(214), I3 =>  inp_feat(206), I4 =>  inp_feat(364), I5 =>  inp_feat(87), I6 =>  inp_feat(90), I7 =>  inp_feat(305)); 
C_49_S_2_L_2_inst : LUT8 generic map(INIT => "1000000010100000111100011010000000100000101000001100000010100000000000001111001000000000000000001000000010000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_2_L_2_out, I0 =>  inp_feat(340), I1 =>  inp_feat(439), I2 =>  inp_feat(435), I3 =>  inp_feat(183), I4 =>  inp_feat(105), I5 =>  inp_feat(74), I6 =>  inp_feat(128), I7 =>  inp_feat(305)); 
C_49_S_2_L_3_inst : LUT8 generic map(INIT => "1111111110001000001101000000000000101001100100000001000000000000000001000000110010001000010000000110000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_2_L_3_out, I0 =>  inp_feat(210), I1 =>  inp_feat(41), I2 =>  inp_feat(161), I3 =>  inp_feat(198), I4 =>  inp_feat(328), I5 =>  inp_feat(364), I6 =>  inp_feat(221), I7 =>  inp_feat(305)); 
C_49_S_2_L_4_inst : LUT8 generic map(INIT => "1010101010101000000000001000000000001000001010101000100011100010101000000000000000000000000000000000100000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_2_L_4_out, I0 =>  inp_feat(230), I1 =>  inp_feat(384), I2 =>  inp_feat(74), I3 =>  inp_feat(80), I4 =>  inp_feat(328), I5 =>  inp_feat(390), I6 =>  inp_feat(227), I7 =>  inp_feat(305)); 
C_49_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000000000000000000000000000000000000010000001111110000010001111100000000010101000000000000000111000000000101010100000001000100010000000000000001000000000000000000100111110001110100010000000000000000000000010100000101000000000") port map( O =>C_49_S_2_L_5_out, I0 =>  inp_feat(473), I1 =>  inp_feat(263), I2 =>  inp_feat(216), I3 =>  inp_feat(106), I4 =>  inp_feat(130), I5 =>  inp_feat(12), I6 =>  inp_feat(323), I7 =>  inp_feat(71)); 
C_49_S_2_L_6_inst : LUT8 generic map(INIT => "0000000110000101000000010000100110110011101010001100001000000000000000000000000000000000100000000000000000000000000000000000000000001000000000010000100000000000100010000000100010000000000000000000000000000000000000000000000011000000000000000000000010000000") port map( O =>C_49_S_2_L_6_out, I0 =>  inp_feat(6), I1 =>  inp_feat(182), I2 =>  inp_feat(451), I3 =>  inp_feat(111), I4 =>  inp_feat(340), I5 =>  inp_feat(290), I6 =>  inp_feat(470), I7 =>  inp_feat(370)); 
C_49_S_2_L_7_inst : LUT8 generic map(INIT => "0010100000100000000000000000000000101011000100000000100000000000000010000000000000000000000000000000000000000000000000000000000011101000000000100010101000000000111011000010011000000101001000001000100000000000000000000000000010000000101000000000000000000000") port map( O =>C_49_S_2_L_7_out, I0 =>  inp_feat(210), I1 =>  inp_feat(259), I2 =>  inp_feat(382), I3 =>  inp_feat(328), I4 =>  inp_feat(470), I5 =>  inp_feat(380), I6 =>  inp_feat(221), I7 =>  inp_feat(95)); 
C_49_S_3_L_0_inst : LUT8 generic map(INIT => "0011010101010000100000000001010001000000000000110100001000000010001111000101110001100001000000101101111100001010011111100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_49_S_3_L_0_out, I0 =>  inp_feat(183), I1 =>  inp_feat(11), I2 =>  inp_feat(362), I3 =>  inp_feat(449), I4 =>  inp_feat(285), I5 =>  inp_feat(54), I6 =>  inp_feat(267), I7 =>  inp_feat(305)); 
C_49_S_3_L_1_inst : LUT8 generic map(INIT => "0010000000000010101100001010000000000000000000000000000000000000100000000000001000001010000000100000000000000000000000000000001010000000001000100110000010100001000000011011101011010000111101001000000000000000000000000010000000000000000000000000000000000000") port map( O =>C_49_S_3_L_1_out, I0 =>  inp_feat(473), I1 =>  inp_feat(87), I2 =>  inp_feat(317), I3 =>  inp_feat(216), I4 =>  inp_feat(267), I5 =>  inp_feat(214), I6 =>  inp_feat(374), I7 =>  inp_feat(160)); 
C_49_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000010000100100000011000100000000000101110100000101000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_3_L_2_out, I0 =>  inp_feat(224), I1 =>  inp_feat(374), I2 =>  inp_feat(76), I3 =>  inp_feat(112), I4 =>  inp_feat(466), I5 =>  inp_feat(381), I6 =>  inp_feat(22), I7 =>  inp_feat(40)); 
C_49_S_3_L_3_inst : LUT8 generic map(INIT => "0000001010000000000000000000000011100010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010111100000000000011000000111000001010000000000000100000000000000000000000000000000000000000000000010000000000000000000000") port map( O =>C_49_S_3_L_3_out, I0 =>  inp_feat(435), I1 =>  inp_feat(460), I2 =>  inp_feat(433), I3 =>  inp_feat(207), I4 =>  inp_feat(46), I5 =>  inp_feat(267), I6 =>  inp_feat(40), I7 =>  inp_feat(365)); 
C_49_S_3_L_4_inst : LUT8 generic map(INIT => "0010000000000100011101010000000000000000000000000000000000000000110110110100010000110001000000000000000000000010001000000000000000000000000000010000000000000000000000000000001000000000000000000000001000000010000000000000000000000000000000000000000000000000") port map( O =>C_49_S_3_L_4_out, I0 =>  inp_feat(480), I1 =>  inp_feat(376), I2 =>  inp_feat(1), I3 =>  inp_feat(282), I4 =>  inp_feat(27), I5 =>  inp_feat(205), I6 =>  inp_feat(5), I7 =>  inp_feat(322)); 
C_49_S_3_L_5_inst : LUT8 generic map(INIT => "1110010010110000110100100100000000000000110000001000000000000000000000000101010000000000000000001100000011000000110000000000000000000001000000010000000000010000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000") port map( O =>C_49_S_3_L_5_out, I0 =>  inp_feat(65), I1 =>  inp_feat(103), I2 =>  inp_feat(378), I3 =>  inp_feat(203), I4 =>  inp_feat(390), I5 =>  inp_feat(504), I6 =>  inp_feat(111), I7 =>  inp_feat(322)); 
C_49_S_3_L_6_inst : LUT8 generic map(INIT => "1000100010101000000000000100101000001000100000000000000000100000000000001100100000000000100000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_3_L_6_out, I0 =>  inp_feat(154), I1 =>  inp_feat(46), I2 =>  inp_feat(329), I3 =>  inp_feat(108), I4 =>  inp_feat(130), I5 =>  inp_feat(143), I6 =>  inp_feat(322), I7 =>  inp_feat(305)); 
C_49_S_3_L_7_inst : LUT8 generic map(INIT => "1111111011100000001000000000000011110011001001010000010000000000110010001111000010010010001100001100001100100001000000000011000000000000000000000000000000000000000000000000000000000000000000001000000001010101000000000000000000000000000100010000000000010001") port map( O =>C_49_S_3_L_7_out, I0 =>  inp_feat(263), I1 =>  inp_feat(103), I2 =>  inp_feat(317), I3 =>  inp_feat(234), I4 =>  inp_feat(130), I5 =>  inp_feat(384), I6 =>  inp_feat(108), I7 =>  inp_feat(322)); 
C_49_S_4_L_0_inst : LUT8 generic map(INIT => "0000110001000000000000000000000000001100000000000000000000000000000011000000000010100000000000000000010000000000000000000000000001000100000000000100010000000000100000000100000000000000000000000100110000000000000000000000000011001100000000000000000000000000") port map( O =>C_49_S_4_L_0_out, I0 =>  inp_feat(71), I1 =>  inp_feat(230), I2 =>  inp_feat(216), I3 =>  inp_feat(46), I4 =>  inp_feat(328), I5 =>  inp_feat(461), I6 =>  inp_feat(160), I7 =>  inp_feat(408)); 
C_49_S_4_L_1_inst : LUT8 generic map(INIT => "0001000000000000000000000000000000000000001100100000000000000000101000001000001000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_4_L_1_out, I0 =>  inp_feat(46), I1 =>  inp_feat(218), I2 =>  inp_feat(40), I3 =>  inp_feat(496), I4 =>  inp_feat(486), I5 =>  inp_feat(340), I6 =>  inp_feat(487), I7 =>  inp_feat(305)); 
C_49_S_4_L_2_inst : LUT8 generic map(INIT => "1010101000000000100000100001101000001111000000000000001100000000000110110000100011111111001011010000000000001100001010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_4_L_2_out, I0 =>  inp_feat(52), I1 =>  inp_feat(120), I2 =>  inp_feat(71), I3 =>  inp_feat(340), I4 =>  inp_feat(62), I5 =>  inp_feat(500), I6 =>  inp_feat(74), I7 =>  inp_feat(305)); 
C_49_S_4_L_3_inst : LUT8 generic map(INIT => "0010000011100000000100010010000000000000010010000000000010000000001011111110000000011010100000000000000011000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000") port map( O =>C_49_S_4_L_3_out, I0 =>  inp_feat(328), I1 =>  inp_feat(316), I2 =>  inp_feat(283), I3 =>  inp_feat(428), I4 =>  inp_feat(29), I5 =>  inp_feat(479), I6 =>  inp_feat(483), I7 =>  inp_feat(151)); 
C_49_S_4_L_4_inst : LUT8 generic map(INIT => "0010011010001101000000000000000001011100100011010000000000000010100000001101011110000000100000000000100011011101000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000") port map( O =>C_49_S_4_L_4_out, I0 =>  inp_feat(7), I1 =>  inp_feat(107), I2 =>  inp_feat(198), I3 =>  inp_feat(183), I4 =>  inp_feat(214), I5 =>  inp_feat(296), I6 =>  inp_feat(80), I7 =>  inp_feat(151)); 
C_49_S_4_L_5_inst : LUT8 generic map(INIT => "0011001000000011000000000000000000010010000000000000000000000000101001110010101000000010000000100110111000000010000000100000101000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000001000000000000000000000000000") port map( O =>C_49_S_4_L_5_out, I0 =>  inp_feat(423), I1 =>  inp_feat(71), I2 =>  inp_feat(387), I3 =>  inp_feat(428), I4 =>  inp_feat(46), I5 =>  inp_feat(130), I6 =>  inp_feat(108), I7 =>  inp_feat(322)); 
C_49_S_4_L_6_inst : LUT8 generic map(INIT => "0010100110000010001010100000100000000000000000000000000000000010001010100000100010101111000000000000000000000010100010000000001000000010000000000100000000000000000000000000000000000000000000000010000000000000001000000001000000000000000000000010000000000001") port map( O =>C_49_S_4_L_6_out, I0 =>  inp_feat(109), I1 =>  inp_feat(80), I2 =>  inp_feat(1), I3 =>  inp_feat(349), I4 =>  inp_feat(316), I5 =>  inp_feat(91), I6 =>  inp_feat(504), I7 =>  inp_feat(227)); 
C_49_S_4_L_7_inst : LUT8 generic map(INIT => "1011101000001111101010000001100000101000000000001010110000100000000010000000000000001000000000100000000000000000001000000000000000010000000000000000110000000000000000000000000000000000000000000000000000000100000000000000010010000000000000000000000000000000") port map( O =>C_49_S_4_L_7_out, I0 =>  inp_feat(451), I1 =>  inp_feat(467), I2 =>  inp_feat(54), I3 =>  inp_feat(15), I4 =>  inp_feat(428), I5 =>  inp_feat(466), I6 =>  inp_feat(79), I7 =>  inp_feat(327)); 
C_50_S_0_L_0_inst : LUT8 generic map(INIT => "1111101111101111111110001111111110001010000011110000000010000111111110000000100001110000001110110000000000000000000000000000000011000000100000101100000000000000000000100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_50_S_0_L_0_out, I0 =>  inp_feat(229), I1 =>  inp_feat(46), I2 =>  inp_feat(40), I3 =>  inp_feat(161), I4 =>  inp_feat(373), I5 =>  inp_feat(332), I6 =>  inp_feat(296), I7 =>  inp_feat(111)); 
C_50_S_0_L_1_inst : LUT8 generic map(INIT => "1110111010100000101000000000100010100100100011000000110000001100011010101000101010101000000010100010110010101110000011001000110000001110100001001000100000000000000010111100110000000100000000000000110010001000100001000000000000000101110011001000010010000110") port map( O =>C_50_S_0_L_1_out, I0 =>  inp_feat(198), I1 =>  inp_feat(183), I2 =>  inp_feat(317), I3 =>  inp_feat(214), I4 =>  inp_feat(216), I5 =>  inp_feat(266), I6 =>  inp_feat(200), I7 =>  inp_feat(71)); 
C_50_S_0_L_2_inst : LUT8 generic map(INIT => "1111111110110000111010000010000000001000000000001010111000000000111111001111010010110000001000000000010000000000001000000000000011010111000000000101100000000000010100000000000001101100001000001101011100000000111111110000000000100011000000001011001100100010") port map( O =>C_50_S_0_L_2_out, I0 =>  inp_feat(493), I1 =>  inp_feat(479), I2 =>  inp_feat(229), I3 =>  inp_feat(267), I4 =>  inp_feat(81), I5 =>  inp_feat(66), I6 =>  inp_feat(40), I7 =>  inp_feat(310)); 
C_50_S_0_L_3_inst : LUT8 generic map(INIT => "0110001011111000000000001010000000111011100000000010000010000000101100001010000000000000100000001111001000000000000000001000000011111010111100001110000011110000100000001100000011000000110000000100000011110000000000001101000000000000010000000000000000000000") port map( O =>C_50_S_0_L_3_out, I0 =>  inp_feat(87), I1 =>  inp_feat(474), I2 =>  inp_feat(74), I3 =>  inp_feat(170), I4 =>  inp_feat(60), I5 =>  inp_feat(436), I6 =>  inp_feat(157), I7 =>  inp_feat(492)); 
C_50_S_0_L_4_inst : LUT8 generic map(INIT => "0010111011111010110111100011000010111000111000000011001000010000111000111110001011100011101000100010001001100010000000000000000000010001000100100000001101000000001100000001000000010011000100000010001100100011000000110000000000100001000000110000001000000000") port map( O =>C_50_S_0_L_4_out, I0 =>  inp_feat(362), I1 =>  inp_feat(364), I2 =>  inp_feat(422), I3 =>  inp_feat(221), I4 =>  inp_feat(355), I5 =>  inp_feat(483), I6 =>  inp_feat(492), I7 =>  inp_feat(408)); 
C_50_S_0_L_5_inst : LUT8 generic map(INIT => "1111110011100000110001001000010010000000110101000100000001000000110011001101110101010100010101001101000011010100000001000100000011111100110011000100100000001100110111011101110101100100000111011100110011001100000001000000100011000000110001000000000000000000") port map( O =>C_50_S_0_L_5_out, I0 =>  inp_feat(435), I1 =>  inp_feat(439), I2 =>  inp_feat(87), I3 =>  inp_feat(479), I4 =>  inp_feat(483), I5 =>  inp_feat(504), I6 =>  inp_feat(448), I7 =>  inp_feat(151)); 
C_50_S_0_L_6_inst : LUT8 generic map(INIT => "1101101010010000110000001110010011000000000000001100000010000000111111101000100011011100111110001001000011100000110011001111000010001000000000000000000010001000101000000000000000000000000000001111000000000000000000001111000011110000100000001100000010100000") port map( O =>C_50_S_0_L_6_out, I0 =>  inp_feat(373), I1 =>  inp_feat(105), I2 =>  inp_feat(183), I3 =>  inp_feat(368), I4 =>  inp_feat(241), I5 =>  inp_feat(74), I6 =>  inp_feat(340), I7 =>  inp_feat(316)); 
C_50_S_0_L_7_inst : LUT8 generic map(INIT => "0101111111000101110111000000000000001100101000000000110000000000010011011111111100000100100000100000010010101000000001000000010011011111110010001100110010000001100010001000100010001100100010001101111010001000110111010000000000001000100000000000111010001000") port map( O =>C_50_S_0_L_7_out, I0 =>  inp_feat(396), I1 =>  inp_feat(439), I2 =>  inp_feat(475), I3 =>  inp_feat(266), I4 =>  inp_feat(87), I5 =>  inp_feat(271), I6 =>  inp_feat(267), I7 =>  inp_feat(151)); 
C_50_S_1_L_0_inst : LUT8 generic map(INIT => "1110110010110000111011110000000010001000101010000100110000000000101001001011100110111111101111010000100010101000000011000000001010000001111000001010111100001000000000001010000000000000000000001101000011010000101101001010001000001100101011100000000011001110") port map( O =>C_50_S_1_L_0_out, I0 =>  inp_feat(373), I1 =>  inp_feat(331), I2 =>  inp_feat(365), I3 =>  inp_feat(220), I4 =>  inp_feat(340), I5 =>  inp_feat(310), I6 =>  inp_feat(200), I7 =>  inp_feat(71)); 
C_50_S_1_L_1_inst : LUT8 generic map(INIT => "0111111111111011110100100111101111101000111010001100000000000000001000001011101000000000001000000110000000100000010000000000000010101000101010001110000010100000101010001010100000000000000000000010000000100000000000000000000010100000001000000000000000000000") port map( O =>C_50_S_1_L_1_out, I0 =>  inp_feat(428), I1 =>  inp_feat(15), I2 =>  inp_feat(158), I3 =>  inp_feat(473), I4 =>  inp_feat(267), I5 =>  inp_feat(151), I6 =>  inp_feat(183), I7 =>  inp_feat(305)); 
C_50_S_1_L_2_inst : LUT8 generic map(INIT => "0010010000000000011011000100010011111110000000000010111000000000101010101000000010101010101010101010101000001000001000100000000011101100000001000100110000001100101100000000000000000000000000001010000010000000000000000000000010100000000000000000000000000000") port map( O =>C_50_S_1_L_2_out, I0 =>  inp_feat(113), I1 =>  inp_feat(387), I2 =>  inp_feat(23), I3 =>  inp_feat(439), I4 =>  inp_feat(436), I5 =>  inp_feat(157), I6 =>  inp_feat(492), I7 =>  inp_feat(305)); 
C_50_S_1_L_3_inst : LUT8 generic map(INIT => "1011001100100011111000001010000111111000110000001110000011010000101110110010001101110010000000111111001000000000001000000000000011000000100000000000000000000000110010001000100000000000000000001010001000000000101010100000101010100010000000000000000000000000") port map( O =>C_50_S_1_L_3_out, I0 =>  inp_feat(87), I1 =>  inp_feat(340), I2 =>  inp_feat(187), I3 =>  inp_feat(439), I4 =>  inp_feat(267), I5 =>  inp_feat(151), I6 =>  inp_feat(221), I7 =>  inp_feat(305)); 
C_50_S_1_L_4_inst : LUT8 generic map(INIT => "1111011111001000111111011101000011110101000000000100000000000000100010001000000001000000000000001111100000000000000000000000000011001100000000001110100010110000000010010000000011000000000000001000100010000000110010000000000000000000000000001000000000000000") port map( O =>C_50_S_1_L_4_out, I0 =>  inp_feat(302), I1 =>  inp_feat(373), I2 =>  inp_feat(1), I3 =>  inp_feat(413), I4 =>  inp_feat(285), I5 =>  inp_feat(54), I6 =>  inp_feat(305), I7 =>  inp_feat(316)); 
C_50_S_1_L_5_inst : LUT8 generic map(INIT => "1111111111111111111111111000111100011001110011111100111001000101100010101010101010000000000000000000001000100000000000000000000010100001001010100000000000001010000000000000000000000000000000001000001000101010100000001000100000000000000000000000000000000000") port map( O =>C_50_S_1_L_5_out, I0 =>  inp_feat(120), I1 =>  inp_feat(7), I2 =>  inp_feat(86), I3 =>  inp_feat(298), I4 =>  inp_feat(198), I5 =>  inp_feat(183), I6 =>  inp_feat(137), I7 =>  inp_feat(60)); 
C_50_S_1_L_6_inst : LUT8 generic map(INIT => "0011110101010011100001110000000011110001001001110000000000000010111101111111000100000100000000001000000110000011000000000000000011101000101010101000010000000000111000001010001000000000001000101100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_50_S_1_L_6_out, I0 =>  inp_feat(109), I1 =>  inp_feat(41), I2 =>  inp_feat(328), I3 =>  inp_feat(407), I4 =>  inp_feat(439), I5 =>  inp_feat(373), I6 =>  inp_feat(111), I7 =>  inp_feat(322)); 
C_50_S_1_L_7_inst : LUT8 generic map(INIT => "1110110111001101110111011111010101100100110101101101010101111100111011001110000011110101000000001100000011100000111101001100000011100000111000000000010100000000010101011101010100000100000000001100110000100000011101010010000000000000000000000011000100000000") port map( O =>C_50_S_1_L_7_out, I0 =>  inp_feat(52), I1 =>  inp_feat(105), I2 =>  inp_feat(152), I3 =>  inp_feat(5), I4 =>  inp_feat(310), I5 =>  inp_feat(201), I6 =>  inp_feat(40), I7 =>  inp_feat(480)); 
C_50_S_2_L_0_inst : LUT8 generic map(INIT => "1011110101111010001111000000000011010011000000000001001100000000111111110111101000011000000000000000000000000000000000000000000011111010000000001111100000000000110010000000000000000000000000000100100000000000111110000000000000001000000000000000000000000000") port map( O =>C_50_S_2_L_0_out, I0 =>  inp_feat(475), I1 =>  inp_feat(396), I2 =>  inp_feat(288), I3 =>  inp_feat(60), I4 =>  inp_feat(135), I5 =>  inp_feat(213), I6 =>  inp_feat(247), I7 =>  inp_feat(305)); 
C_50_S_2_L_1_inst : LUT8 generic map(INIT => "0100100011001100101010100000000011101101010011001110111000000100100000011000110000000000000000000000111000001100000000000000010011101010110010101110101010000000101010101000101000001010000000000000101011001110000000000000000010001010110011100000000000000000") port map( O =>C_50_S_2_L_1_out, I0 =>  inp_feat(33), I1 =>  inp_feat(87), I2 =>  inp_feat(15), I3 =>  inp_feat(143), I4 =>  inp_feat(205), I5 =>  inp_feat(473), I6 =>  inp_feat(203), I7 =>  inp_feat(492)); 
C_50_S_2_L_2_inst : LUT8 generic map(INIT => "0100001000000000101110010000001010011010001100001111001000000010101000000011000010000000000000001010000000000000000000000000000011111100111100001111110110100000101100101111101011111010001010101111000011110000000000000000000011000000011100000000000000000000") port map( O =>C_50_S_2_L_2_out, I0 =>  inp_feat(353), I1 =>  inp_feat(362), I2 =>  inp_feat(74), I3 =>  inp_feat(87), I4 =>  inp_feat(340), I5 =>  inp_feat(390), I6 =>  inp_feat(486), I7 =>  inp_feat(328)); 
C_50_S_2_L_3_inst : LUT8 generic map(INIT => "0111010011101000000000000010000010100010001000101010000000000000101110110111000000100001000000000010001010100010100000000000000011100110110101000100000000000000111001001111110111000000010000000000000000000000000000000000000011011000111111011100000000000000") port map( O =>C_50_S_2_L_3_out, I0 =>  inp_feat(422), I1 =>  inp_feat(362), I2 =>  inp_feat(483), I3 =>  inp_feat(469), I4 =>  inp_feat(267), I5 =>  inp_feat(40), I6 =>  inp_feat(428), I7 =>  inp_feat(492)); 
C_50_S_2_L_4_inst : LUT8 generic map(INIT => "1111101011111010111111111110001110000000000000000010001000100000100000000001101000101010111100010000000000000000100000100000000011111110111111001110111011111100011000001101110011100010110011000010000011111010101000101110100010001000100010001010001010001000") port map( O =>C_50_S_2_L_4_out, I0 =>  inp_feat(120), I1 =>  inp_feat(310), I2 =>  inp_feat(373), I3 =>  inp_feat(5), I4 =>  inp_feat(340), I5 =>  inp_feat(480), I6 =>  inp_feat(105), I7 =>  inp_feat(221)); 
C_50_S_2_L_5_inst : LUT8 generic map(INIT => "1110111011101110111010101010111111001100101011100100100010000101110000000010000010001000100010001100100000000000110010000000000011111010111011100010101010100000111010111010101100001110100010000100100000000000000010000000000000001000000000001100101000000000") port map( O =>C_50_S_2_L_5_out, I0 =>  inp_feat(436), I1 =>  inp_feat(452), I2 =>  inp_feat(15), I3 =>  inp_feat(218), I4 =>  inp_feat(233), I5 =>  inp_feat(408), I6 =>  inp_feat(437), I7 =>  inp_feat(149)); 
C_50_S_2_L_6_inst : LUT8 generic map(INIT => "1100100011101010100010001111110011000101111000001000000010101010110010001110001000001000111000101000110001101010000010001100100011000000011000001010100011100010000100111010001010001010000000000000000000000010000010000000000000000000000100010000101000111000") port map( O =>C_50_S_2_L_6_out, I0 =>  inp_feat(480), I1 =>  inp_feat(138), I2 =>  inp_feat(367), I3 =>  inp_feat(180), I4 =>  inp_feat(331), I5 =>  inp_feat(483), I6 =>  inp_feat(161), I7 =>  inp_feat(390)); 
C_50_S_2_L_7_inst : LUT8 generic map(INIT => "1111111110111111011000001010000010001100101110010000010000000000111000001010111000100010101001001000000010001000000000000000000011110111011101111101010000000000011101011111010101010100010101001110010011101100010000000100010010010100011111100000000000000000") port map( O =>C_50_S_2_L_7_out, I0 =>  inp_feat(34), I1 =>  inp_feat(178), I2 =>  inp_feat(297), I3 =>  inp_feat(418), I4 =>  inp_feat(74), I5 =>  inp_feat(11), I6 =>  inp_feat(267), I7 =>  inp_feat(151)); 
C_50_S_3_L_0_inst : LUT8 generic map(INIT => "0111011001010000111100001101000010110011101100101111000010000000110011110000000111000111110000110000000000000000111111111100000111101010000000001100000010000000101010101010101000000000000000000000000000000000110000000000000000000000000000000000000000000000") port map( O =>C_50_S_3_L_0_out, I0 =>  inp_feat(15), I1 =>  inp_feat(100), I2 =>  inp_feat(232), I3 =>  inp_feat(267), I4 =>  inp_feat(40), I5 =>  inp_feat(428), I6 =>  inp_feat(492), I7 =>  inp_feat(151)); 
C_50_S_3_L_1_inst : LUT8 generic map(INIT => "0110100011101010100010001000000011110000110000001010000011000000101010101110000000000000100000001101000011110000010000000000000010011000010010100000100000001000111110101111101001001000110010000000000000000000000000000000000010111010111110100000000000001000") port map( O =>C_50_S_3_L_1_out, I0 =>  inp_feat(90), I1 =>  inp_feat(285), I2 =>  inp_feat(422), I3 =>  inp_feat(329), I4 =>  inp_feat(342), I5 =>  inp_feat(40), I6 =>  inp_feat(428), I7 =>  inp_feat(492)); 
C_50_S_3_L_2_inst : LUT8 generic map(INIT => "0111100110101000111010010000000010101100101010101110000000000000110011101000100001001100001010101100111000001000011000000000000011111111000010101000101000101010001000100000001000100010000000100110111100000010001010100010101000100010000000100000000000000000") port map( O =>C_50_S_3_L_2_out, I0 =>  inp_feat(287), I1 =>  inp_feat(310), I2 =>  inp_feat(15), I3 =>  inp_feat(229), I4 =>  inp_feat(428), I5 =>  inp_feat(436), I6 =>  inp_feat(157), I7 =>  inp_feat(492)); 
C_50_S_3_L_3_inst : LUT8 generic map(INIT => "1011111110000000111111011000100010100011101010101000111100001110000101110000110010001111100010000001010100000000000001010000000010110101000001000011110000001000101001101010111000000110000011100000100100001100000000000000110000000100000001000000010000001100") port map( O =>C_50_S_3_L_3_out, I0 =>  inp_feat(88), I1 =>  inp_feat(156), I2 =>  inp_feat(328), I3 =>  inp_feat(183), I4 =>  inp_feat(298), I5 =>  inp_feat(216), I6 =>  inp_feat(267), I7 =>  inp_feat(151)); 
C_50_S_3_L_4_inst : LUT8 generic map(INIT => "1110101010000000110011111100000011001010100000001100101000001000111010001010100011101010100010000010100000000000000010001000100011001100110010001100000011000100110011011000000011011100110011011010001001000110010010101100000000011000100000000000000010001010") port map( O =>C_50_S_3_L_4_out, I0 =>  inp_feat(368), I1 =>  inp_feat(183), I2 =>  inp_feat(351), I3 =>  inp_feat(365), I4 =>  inp_feat(340), I5 =>  inp_feat(238), I6 =>  inp_feat(290), I7 =>  inp_feat(210)); 
C_50_S_3_L_5_inst : LUT8 generic map(INIT => "0011101011111000000000001000000011111110111110100000001010001000011011101000101000001100000010000000101000001010000010000000100000000000000000000000000000000000101010100000101000001000100010100110101000000000000000000000000000001010000010100000100000001000") port map( O =>C_50_S_3_L_5_out, I0 =>  inp_feat(90), I1 =>  inp_feat(157), I2 =>  inp_feat(46), I3 =>  inp_feat(465), I4 =>  inp_feat(439), I5 =>  inp_feat(191), I6 =>  inp_feat(221), I7 =>  inp_feat(294)); 
C_50_S_3_L_6_inst : LUT8 generic map(INIT => "0101011001110000110011011100100110110011001100011011111100010111000001000110101100001100000011001010111100011111100011110010111100000000000000000100100001000100000000001000001011000101000101010000100000000100000011000000010000001000100000000000100010000000") port map( O =>C_50_S_3_L_6_out, I0 =>  inp_feat(164), I1 =>  inp_feat(220), I2 =>  inp_feat(178), I3 =>  inp_feat(161), I4 =>  inp_feat(470), I5 =>  inp_feat(41), I6 =>  inp_feat(221), I7 =>  inp_feat(294)); 
C_50_S_3_L_7_inst : LUT8 generic map(INIT => "1101111010001111010001101010001011111011010011001101110101101111111111110000010001100101000000001011111110001100111111011000110010010000000011001100010100000000010001101000000010110011011110001111111100000000010101010000000011011100101001011111111101001001") port map( O =>C_50_S_3_L_7_out, I0 =>  inp_feat(41), I1 =>  inp_feat(53), I2 =>  inp_feat(221), I3 =>  inp_feat(42), I4 =>  inp_feat(83), I5 =>  inp_feat(5), I6 =>  inp_feat(52), I7 =>  inp_feat(290)); 
C_50_S_4_L_0_inst : LUT8 generic map(INIT => "0111110011110000100100001001000011111101011101011101010101010000110011001000000001110001100000001010100000000000100010000000000001011000011100001111000000000000011000000101010010000000010100001100000010000000010101000000000000000000000000000000000000000000") port map( O =>C_50_S_4_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(494), I2 =>  inp_feat(439), I3 =>  inp_feat(469), I4 =>  inp_feat(428), I5 =>  inp_feat(492), I6 =>  inp_feat(149), I7 =>  inp_feat(483)); 
C_50_S_4_L_1_inst : LUT8 generic map(INIT => "1100111011000000100000001000000011011100110010001000100000001000110010101101010000001000111101111101110001011100000010001101111100001010000000000000100000000000110101000000000000001000000000000000101000000000000000000000000000000000000000000000100000000000") port map( O =>C_50_S_4_L_1_out, I0 =>  inp_feat(40), I1 =>  inp_feat(439), I2 =>  inp_feat(172), I3 =>  inp_feat(191), I4 =>  inp_feat(294), I5 =>  inp_feat(221), I6 =>  inp_feat(414), I7 =>  inp_feat(149)); 
C_50_S_4_L_2_inst : LUT8 generic map(INIT => "1110110110110100111111011111110011000000000000001001110111101000110111010001010010001101000111001011101100000010010111000110100011000100110001001101110100001000010000000000000000000000000000000000110100000101000001000001110000000000000000000000000000000000") port map( O =>C_50_S_4_L_2_out, I0 =>  inp_feat(142), I1 =>  inp_feat(74), I2 =>  inp_feat(247), I3 =>  inp_feat(373), I4 =>  inp_feat(485), I5 =>  inp_feat(1), I6 =>  inp_feat(316), I7 =>  inp_feat(105)); 
C_50_S_4_L_3_inst : LUT8 generic map(INIT => "1110111111000000111111111100000011111111110000001110101111000000000011000000000010100010010000001000000101000000010000011100000000001100110010001111101011000000101011111100000011001000110000000000100001000000000000000000000001010000100000001100000011000000") port map( O =>C_50_S_4_L_3_out, I0 =>  inp_feat(413), I1 =>  inp_feat(15), I2 =>  inp_feat(212), I3 =>  inp_feat(498), I4 =>  inp_feat(221), I5 =>  inp_feat(227), I6 =>  inp_feat(306), I7 =>  inp_feat(71)); 
C_50_S_4_L_4_inst : LUT8 generic map(INIT => "0001101110100010101110110011001000100000000000001010001000110000110010100000000111101010001100000000000000000000001000000011000010101111000000001010001010100001101000100000000010000010000000000010101100100010001000110010000000100010000000000010001100000000") port map( O =>C_50_S_4_L_4_out, I0 =>  inp_feat(439), I1 =>  inp_feat(84), I2 =>  inp_feat(135), I3 =>  inp_feat(281), I4 =>  inp_feat(298), I5 =>  inp_feat(271), I6 =>  inp_feat(267), I7 =>  inp_feat(151)); 
C_50_S_4_L_5_inst : LUT8 generic map(INIT => "1111111011111000011101001111110110111110001000000000000000000000011011001111101001000101111100101100010000000000000000000000000011111000100010001000000010001010111100000000000000000010000000101010000000000000000000000000001000100000000000000000000000000000") port map( O =>C_50_S_4_L_5_out, I0 =>  inp_feat(475), I1 =>  inp_feat(100), I2 =>  inp_feat(157), I3 =>  inp_feat(46), I4 =>  inp_feat(218), I5 =>  inp_feat(347), I6 =>  inp_feat(398), I7 =>  inp_feat(470)); 
C_50_S_4_L_6_inst : LUT8 generic map(INIT => "1000110011001000011001111111101101101110010000000000000000000000101110111100010010000011110100111010101000000000000000000000000011101000100010000010000010001100111000000000000000000001000000011010000000000000000000000000000100000000000000000000000000000000") port map( O =>C_50_S_4_L_6_out, I0 =>  inp_feat(23), I1 =>  inp_feat(236), I2 =>  inp_feat(157), I3 =>  inp_feat(46), I4 =>  inp_feat(218), I5 =>  inp_feat(347), I6 =>  inp_feat(398), I7 =>  inp_feat(470)); 
C_50_S_4_L_7_inst : LUT8 generic map(INIT => "1110101110100110111100001000000011100101000000001111000011000000111110110100111111110101110001001101000111001000111100001100100010111010001000101010000000100000111000100010001011110000001000001111101111001110111101001100000011110101101100001110000011000000") port map( O =>C_50_S_4_L_7_out, I0 =>  inp_feat(420), I1 =>  inp_feat(328), I2 =>  inp_feat(448), I3 =>  inp_feat(74), I4 =>  inp_feat(164), I5 =>  inp_feat(290), I6 =>  inp_feat(52), I7 =>  inp_feat(71)); 
C_51_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000001110000000000000000000000000000001100000000000100010001010100010111000000000000000000000000000000000000000000000000000000001000000100000000000000001010000010000000000000000000000000000000000100010000000000000000") port map( O =>C_51_S_0_L_0_out, I0 =>  inp_feat(87), I1 =>  inp_feat(33), I2 =>  inp_feat(216), I3 =>  inp_feat(1), I4 =>  inp_feat(266), I5 =>  inp_feat(267), I6 =>  inp_feat(4), I7 =>  inp_feat(368)); 
C_51_S_0_L_1_inst : LUT8 generic map(INIT => "0110000001100101000100000010000000000000000000000000000000000000000010000100010001000000000000000000000000000000000000000000000010100010111110100000011010000010000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_51_S_0_L_1_out, I0 =>  inp_feat(204), I1 =>  inp_feat(267), I2 =>  inp_feat(9), I3 =>  inp_feat(54), I4 =>  inp_feat(340), I5 =>  inp_feat(12), I6 =>  inp_feat(475), I7 =>  inp_feat(155)); 
C_51_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000111000000000000010010000000000000000011000001000101000100000000001000010000000000000000000000000010000000000000011110000000000000100010100000010") port map( O =>C_51_S_0_L_2_out, I0 =>  inp_feat(267), I1 =>  inp_feat(86), I2 =>  inp_feat(157), I3 =>  inp_feat(239), I4 =>  inp_feat(27), I5 =>  inp_feat(87), I6 =>  inp_feat(296), I7 =>  inp_feat(4)); 
C_51_S_0_L_3_inst : LUT8 generic map(INIT => "0110000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001110111000011010000011100000101000000000000000000000000000000000101111100001111001010110000001000000000000000000000000000000000") port map( O =>C_51_S_0_L_3_out, I0 =>  inp_feat(66), I1 =>  inp_feat(7), I2 =>  inp_feat(247), I3 =>  inp_feat(152), I4 =>  inp_feat(223), I5 =>  inp_feat(40), I6 =>  inp_feat(402), I7 =>  inp_feat(4)); 
C_51_S_0_L_4_inst : LUT8 generic map(INIT => "0000100000000000000000000000000000001000000000000010000000000000000000000000000001101000000000000100100000000000000011100000000000000000000000000000000000000000100000000000000010101010000001011000011100000001000111010001100110000000000000001101111000000000") port map( O =>C_51_S_0_L_4_out, I0 =>  inp_feat(493), I1 =>  inp_feat(460), I2 =>  inp_feat(87), I3 =>  inp_feat(435), I4 =>  inp_feat(439), I5 =>  inp_feat(420), I6 =>  inp_feat(71), I7 =>  inp_feat(4)); 
C_51_S_0_L_5_inst : LUT8 generic map(INIT => "0000000110000000000000000000000000000000101010000000100000001000000000000000000000000000000000000000000000000000000000000000000000010001001000100011001100010011011001111010101100010001000111010000001000000000000000000000000100000110000011100000000000000000") port map( O =>C_51_S_0_L_5_out, I0 =>  inp_feat(15), I1 =>  inp_feat(54), I2 =>  inp_feat(387), I3 =>  inp_feat(365), I4 =>  inp_feat(329), I5 =>  inp_feat(108), I6 =>  inp_feat(143), I7 =>  inp_feat(333)); 
C_51_S_0_L_6_inst : LUT8 generic map(INIT => "0010101000000011110100100010001000000000000000001000100000000000111000000000000000100000101010100000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000010000000") port map( O =>C_51_S_0_L_6_out, I0 =>  inp_feat(186), I1 =>  inp_feat(201), I2 =>  inp_feat(207), I3 =>  inp_feat(291), I4 =>  inp_feat(183), I5 =>  inp_feat(481), I6 =>  inp_feat(74), I7 =>  inp_feat(151)); 
C_51_S_0_L_7_inst : LUT8 generic map(INIT => "0110001101010101001000001000001100000000101001110101001000110010000000000001000000000000000000000001100000011010001110000001001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000001000100010001000100010") port map( O =>C_51_S_0_L_7_out, I0 =>  inp_feat(238), I1 =>  inp_feat(286), I2 =>  inp_feat(82), I3 =>  inp_feat(365), I4 =>  inp_feat(65), I5 =>  inp_feat(105), I6 =>  inp_feat(35), I7 =>  inp_feat(492)); 
C_51_S_1_L_0_inst : LUT8 generic map(INIT => "0000111010001100000010000010100001010011000000000000000000101010000000000000000000001001001010000101100000000010000000101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000") port map( O =>C_51_S_1_L_0_out, I0 =>  inp_feat(362), I1 =>  inp_feat(108), I2 =>  inp_feat(183), I3 =>  inp_feat(439), I4 =>  inp_feat(291), I5 =>  inp_feat(54), I6 =>  inp_feat(285), I7 =>  inp_feat(492)); 
C_51_S_1_L_1_inst : LUT8 generic map(INIT => "0000000001000100000000000000000000000100000010000000000001000000000000000000000000000000000000000000000000000000000000000000000010100100000111011000010010000000000011001100110000000000000000000000000000000000000000000000000000000000000011010000000000000000") port map( O =>C_51_S_1_L_1_out, I0 =>  inp_feat(195), I1 =>  inp_feat(170), I2 =>  inp_feat(333), I3 =>  inp_feat(201), I4 =>  inp_feat(380), I5 =>  inp_feat(332), I6 =>  inp_feat(143), I7 =>  inp_feat(4)); 
C_51_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000010001001101010100000000000000001000101000000000000000000000000011110000111001101000000000000000000001010000000000000000000000001111110111010000000000000000000000001000000000000000000000000000") port map( O =>C_51_S_1_L_2_out, I0 =>  inp_feat(373), I1 =>  inp_feat(340), I2 =>  inp_feat(221), I3 =>  inp_feat(201), I4 =>  inp_feat(132), I5 =>  inp_feat(249), I6 =>  inp_feat(365), I7 =>  inp_feat(138)); 
C_51_S_1_L_3_inst : LUT8 generic map(INIT => "0000010000000000000001000000000011010100010011000000000010000000010001000000100000000100000010101000101000000000000000001000000001000100000000000000000000000000110011001000000010001000000000000000000000000000000010000000000000000000000000001000100000000000") port map( O =>C_51_S_1_L_3_out, I0 =>  inp_feat(296), I1 =>  inp_feat(435), I2 =>  inp_feat(477), I3 =>  inp_feat(67), I4 =>  inp_feat(362), I5 =>  inp_feat(483), I6 =>  inp_feat(62), I7 =>  inp_feat(160)); 
C_51_S_1_L_4_inst : LUT8 generic map(INIT => "0000010000000000000000110000000000000000000000000000000000000000000011000000000001001001000000000000100010000000000000000000000010001001000000000000010000000000100000101000000000101010000000000000000010000000000010001000000010001000100000000000000010000000") port map( O =>C_51_S_1_L_4_out, I0 =>  inp_feat(360), I1 =>  inp_feat(211), I2 =>  inp_feat(71), I3 =>  inp_feat(305), I4 =>  inp_feat(7), I5 =>  inp_feat(158), I6 =>  inp_feat(402), I7 =>  inp_feat(4)); 
C_51_S_1_L_5_inst : LUT8 generic map(INIT => "1000110011001000100000001000000000100010000001001000000000000000000010000011100010111011001000100000000000110000100000000000001100000000000000000000000000000000000000000000000000000000000000000000000000110010000000100000000000000000000000000000000000000000") port map( O =>C_51_S_1_L_5_out, I0 =>  inp_feat(317), I1 =>  inp_feat(222), I2 =>  inp_feat(267), I3 =>  inp_feat(216), I4 =>  inp_feat(9), I5 =>  inp_feat(340), I6 =>  inp_feat(1), I7 =>  inp_feat(12)); 
C_51_S_1_L_6_inst : LUT8 generic map(INIT => "0000001000000000000000000000000000000000000000000000000000000000000010100100000000000010000000000000000000000000000000000000000010000010010000101010101010001010000010000100000000000000100000100000001011000000000000101100000000000000000000000000000000000000") port map( O =>C_51_S_1_L_6_out, I0 =>  inp_feat(322), I1 =>  inp_feat(296), I2 =>  inp_feat(480), I3 =>  inp_feat(247), I4 =>  inp_feat(7), I5 =>  inp_feat(228), I6 =>  inp_feat(402), I7 =>  inp_feat(4)); 
C_51_S_1_L_7_inst : LUT8 generic map(INIT => "0000010010000100000000000010100001000000100000001000000011000000000000000000000000000000000000000000000000000000000000000000000011000100100001000000000010000000100000001100100000001100111010110000000000000000000000001000010000000000010001011000000001001101") port map( O =>C_51_S_1_L_7_out, I0 =>  inp_feat(271), I1 =>  inp_feat(435), I2 =>  inp_feat(107), I3 =>  inp_feat(373), I4 =>  inp_feat(303), I5 =>  inp_feat(504), I6 =>  inp_feat(151), I7 =>  inp_feat(120)); 
C_51_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000100010000000000000000000000000000000000000000000001000001010000010001000100010000000000000000000000000000000000010100010000010001001110010110000000000000000000000000000001000000000000010100000100000001000000000000000000000000000000000000000") port map( O =>C_51_S_2_L_0_out, I0 =>  inp_feat(107), I1 =>  inp_feat(222), I2 =>  inp_feat(220), I3 =>  inp_feat(11), I4 =>  inp_feat(183), I5 =>  inp_feat(12), I6 =>  inp_feat(229), I7 =>  inp_feat(38)); 
C_51_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000100000000000000000000000000000000000000000000000000000000100000011000000010000000000000000000000000000000000000000000000010000000100000011001000000000001000000000000000001000000100110001000100010000001100000000000100000000000000000000000000") port map( O =>C_51_S_2_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(435), I2 =>  inp_feat(318), I3 =>  inp_feat(260), I4 =>  inp_feat(428), I5 =>  inp_feat(492), I6 =>  inp_feat(90), I7 =>  inp_feat(4)); 
C_51_S_2_L_2_inst : LUT8 generic map(INIT => "0001000000110000000000000000000000000000001000000000000000000000000000000011000000000000000100000000000000001000000000000000000000000010001000001010000000000000110100000000000000000000000000001000001100001101000000010010110111011101000110000001101100011111") port map( O =>C_51_S_2_L_2_out, I0 =>  inp_feat(385), I1 =>  inp_feat(66), I2 =>  inp_feat(247), I3 =>  inp_feat(402), I4 =>  inp_feat(7), I5 =>  inp_feat(138), I6 =>  inp_feat(331), I7 =>  inp_feat(4)); 
C_51_S_2_L_3_inst : LUT8 generic map(INIT => "0000000010000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000111010001101100010111110000110000000000010100000110110000000000010001000110000000000100000000000001000000000000000000000") port map( O =>C_51_S_2_L_3_out, I0 =>  inp_feat(9), I1 =>  inp_feat(511), I2 =>  inp_feat(317), I3 =>  inp_feat(90), I4 =>  inp_feat(103), I5 =>  inp_feat(12), I6 =>  inp_feat(340), I7 =>  inp_feat(4)); 
C_51_S_2_L_4_inst : LUT8 generic map(INIT => "0000001000000000000000000000000000000000000000000000000000000000000000110000000000000010000000000001001000000000000000000000000000000011000000010001000100000110101100110000000000000011000101010010001100000000000000100000000000110001000000000111101000000000") port map( O =>C_51_S_2_L_4_out, I0 =>  inp_feat(158), I1 =>  inp_feat(45), I2 =>  inp_feat(66), I3 =>  inp_feat(228), I4 =>  inp_feat(7), I5 =>  inp_feat(138), I6 =>  inp_feat(402), I7 =>  inp_feat(4)); 
C_51_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000110000000000000000000000000000000000000000011000000001000010100000000000000000000000000000000000000000000000101000100010000010001100000000000000000000000000000001000000001100101000001000101000110000001110000000000000000000000100000001") port map( O =>C_51_S_2_L_5_out, I0 =>  inp_feat(358), I1 =>  inp_feat(420), I2 =>  inp_feat(247), I3 =>  inp_feat(228), I4 =>  inp_feat(260), I5 =>  inp_feat(99), I6 =>  inp_feat(71), I7 =>  inp_feat(4)); 
C_51_S_2_L_6_inst : LUT8 generic map(INIT => "1100110011100000101001001000001000000000001000000010000011100010000010100000100000001000001000000000000000110000000010001111100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100011110000") port map( O =>C_51_S_2_L_6_out, I0 =>  inp_feat(111), I1 =>  inp_feat(31), I2 =>  inp_feat(364), I3 =>  inp_feat(267), I4 =>  inp_feat(87), I5 =>  inp_feat(296), I6 =>  inp_feat(260), I7 =>  inp_feat(143)); 
C_51_S_2_L_7_inst : LUT8 generic map(INIT => "0100100000001000000000001010000000001000000000000000000000000000110101001100110001010000010101001101010101010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100010001000000010000000000000000000000") port map( O =>C_51_S_2_L_7_out, I0 =>  inp_feat(49), I1 =>  inp_feat(473), I2 =>  inp_feat(340), I3 =>  inp_feat(90), I4 =>  inp_feat(64), I5 =>  inp_feat(317), I6 =>  inp_feat(1), I7 =>  inp_feat(12)); 
C_51_S_3_L_0_inst : LUT8 generic map(INIT => "0000001000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010110101110000001010000000000000100000001000010010000000001000000000010011001000001010000000000000000000010000000000000000") port map( O =>C_51_S_3_L_0_out, I0 =>  inp_feat(222), I1 =>  inp_feat(387), I2 =>  inp_feat(452), I3 =>  inp_feat(365), I4 =>  inp_feat(163), I5 =>  inp_feat(143), I6 =>  inp_feat(340), I7 =>  inp_feat(4)); 
C_51_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000010000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000001000110001000000000000000000000100000000000000000000000000000000101111101011101111011110000000000000000000000000000100000000000") port map( O =>C_51_S_3_L_1_out, I0 =>  inp_feat(66), I1 =>  inp_feat(234), I2 =>  inp_feat(105), I3 =>  inp_feat(228), I4 =>  inp_feat(402), I5 =>  inp_feat(396), I6 =>  inp_feat(27), I7 =>  inp_feat(4)); 
C_51_S_3_L_2_inst : LUT8 generic map(INIT => "0000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000011100101000000000000000100000001000000000000000000000000000000010000000000000000000000011000000100000000000000000000000") port map( O =>C_51_S_3_L_2_out, I0 =>  inp_feat(239), I1 =>  inp_feat(154), I2 =>  inp_feat(12), I3 =>  inp_feat(90), I4 =>  inp_feat(107), I5 =>  inp_feat(332), I6 =>  inp_feat(143), I7 =>  inp_feat(4)); 
C_51_S_3_L_3_inst : LUT8 generic map(INIT => "0001000000000000000100000000000000000000000000000000000000000000100000000000000010010000110000000000000000000000000000000000000001011000000000000000000000000000100000000000000000000000000000000111001000010001000100000111000100000000000000000000000000000000") port map( O =>C_51_S_3_L_3_out, I0 =>  inp_feat(45), I1 =>  inp_feat(66), I2 =>  inp_feat(152), I3 =>  inp_feat(170), I4 =>  inp_feat(402), I5 =>  inp_feat(396), I6 =>  inp_feat(27), I7 =>  inp_feat(4)); 
C_51_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000100000000000000000000000000000000000000000000001101010000000010010000000000000000000000000000000000010000000110000000000000000000000000000000000000000000000000000000000010011001000100010000000100000000000000000000000000000000000") port map( O =>C_51_S_3_L_4_out, I0 =>  inp_feat(227), I1 =>  inp_feat(425), I2 =>  inp_feat(466), I3 =>  inp_feat(71), I4 =>  inp_feat(402), I5 =>  inp_feat(396), I6 =>  inp_feat(27), I7 =>  inp_feat(4)); 
C_51_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000100000001000000010000000000000000000000000000000000000010001000000000000110000001000000000000000000000000000000000000001110000011000000000000000000000000100001010000000000000000000000010001000100010001100000010000000000000000000000000000000100000") port map( O =>C_51_S_3_L_5_out, I0 =>  inp_feat(271), I1 =>  inp_feat(439), I2 =>  inp_feat(228), I3 =>  inp_feat(460), I4 =>  inp_feat(402), I5 =>  inp_feat(396), I6 =>  inp_feat(27), I7 =>  inp_feat(4)); 
C_51_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100011010000100100000000000000000000000000000000000000000000000010000000001010100000000000000010010001000000100100001100110011001000101000001000000000000000000000001000000000000000100000000000") port map( O =>C_51_S_3_L_6_out, I0 =>  inp_feat(475), I1 =>  inp_feat(227), I2 =>  inp_feat(201), I3 =>  inp_feat(353), I4 =>  inp_feat(239), I5 =>  inp_feat(152), I6 =>  inp_feat(27), I7 =>  inp_feat(4)); 
C_51_S_3_L_7_inst : LUT8 generic map(INIT => "0010110000001000101010000000000100001100000000000000000000000011100011000000100010001010110010111010110010001000000000010000111100000000000000000000000000000000000010000000001000000000000000000000000010000000000000000000000000000010000000000000000100000011") port map( O =>C_51_S_3_L_7_out, I0 =>  inp_feat(340), I1 =>  inp_feat(107), I2 =>  inp_feat(373), I3 =>  inp_feat(418), I4 =>  inp_feat(507), I5 =>  inp_feat(198), I6 =>  inp_feat(504), I7 =>  inp_feat(151)); 
C_51_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000010000000000000001000100000001000000000000000000000000000000000011001101100000001000000000000000000001000000010000000100000000000111010000110101010000010101010100000100000001000000000000000000") port map( O =>C_51_S_4_L_0_out, I0 =>  inp_feat(413), I1 =>  inp_feat(339), I2 =>  inp_feat(182), I3 =>  inp_feat(82), I4 =>  inp_feat(52), I5 =>  inp_feat(456), I6 =>  inp_feat(295), I7 =>  inp_feat(160)); 
C_51_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000110001000000000011000000000000000000000000000000000000000000000000011000111010100001000001000000000000000000000000000100000000000100001000101011110111110000000000000010001000100100010001000000") port map( O =>C_51_S_4_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(477), I2 =>  inp_feat(290), I3 =>  inp_feat(336), I4 =>  inp_feat(260), I5 =>  inp_feat(99), I6 =>  inp_feat(71), I7 =>  inp_feat(4)); 
C_51_S_4_L_2_inst : LUT8 generic map(INIT => "1000000101010101000000000000000000010000000000010000000000000000110111110000000000000100000000001101000010000000010000000000000000000001000100010000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000") port map( O =>C_51_S_4_L_2_out, I0 =>  inp_feat(307), I1 =>  inp_feat(431), I2 =>  inp_feat(291), I3 =>  inp_feat(222), I4 =>  inp_feat(151), I5 =>  inp_feat(107), I6 =>  inp_feat(183), I7 =>  inp_feat(143)); 
C_51_S_4_L_3_inst : LUT8 generic map(INIT => "0010101000001011000000000000000000000010101000000000000000000000001110001010101100000000001010000010101010101111000000000010001100000010000000110000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000") port map( O =>C_51_S_4_L_3_out, I0 =>  inp_feat(435), I1 =>  inp_feat(7), I2 =>  inp_feat(297), I3 =>  inp_feat(87), I4 =>  inp_feat(151), I5 =>  inp_feat(107), I6 =>  inp_feat(183), I7 =>  inp_feat(143)); 
C_51_S_4_L_4_inst : LUT8 generic map(INIT => "1001000010010000000000000000000000000000001010100000000000000000010100001111111100000000001111000101000011010101000000000001000000000000000000000000000000000000000000000010000000000000000000000000000001110010000000000000000000000000000000000000000000000000") port map( O =>C_51_S_4_L_4_out, I0 =>  inp_feat(285), I1 =>  inp_feat(263), I2 =>  inp_feat(317), I3 =>  inp_feat(33), I4 =>  inp_feat(12), I5 =>  inp_feat(64), I6 =>  inp_feat(54), I7 =>  inp_feat(143)); 
C_51_S_4_L_5_inst : LUT8 generic map(INIT => "0000100001000100000000000000000000000000000000001000010000100000000011000100010011000000010001100000000000000100000000100010011000000000000000000000000000000000100010001000100000001000000011000000100000000100000010101010001000000000000001000000010000000100") port map( O =>C_51_S_4_L_5_out, I0 =>  inp_feat(54), I1 =>  inp_feat(107), I2 =>  inp_feat(267), I3 =>  inp_feat(87), I4 =>  inp_feat(88), I5 =>  inp_feat(121), I6 =>  inp_feat(183), I7 =>  inp_feat(303)); 
C_51_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000100011011101000001010000010000001001000001000000000000000000000000000000000000001111010000000000101000000000000000000000001000000010011100110001000000000000000000000000010100000000000000000000000000000000001000000000000000000000000000000000") port map( O =>C_51_S_4_L_6_out, I0 =>  inp_feat(267), I1 =>  inp_feat(373), I2 =>  inp_feat(107), I3 =>  inp_feat(439), I4 =>  inp_feat(71), I5 =>  inp_feat(38), I6 =>  inp_feat(139), I7 =>  inp_feat(303)); 
C_51_S_4_L_7_inst : LUT8 generic map(INIT => "0001001101010101100010101111000100010001000001000000000011011100000000010000000000100110000000010001000000000000000101000101010000011100000000001110001101010100010110100000000010000011000100000000000000000000011111110101010000000011000000000000101100001000") port map( O =>C_51_S_4_L_7_out, I0 =>  inp_feat(71), I1 =>  inp_feat(201), I2 =>  inp_feat(247), I3 =>  inp_feat(152), I4 =>  inp_feat(390), I5 =>  inp_feat(331), I6 =>  inp_feat(83), I7 =>  inp_feat(42)); 
C_52_S_0_L_0_inst : LUT8 generic map(INIT => "1111110010101000111011001000000011001000110000001111101100110110101010000000000010101100000000001000100010000000000000000000000011110000010100001000000010000000110110000001000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_52_S_0_L_0_out, I0 =>  inp_feat(267), I1 =>  inp_feat(173), I2 =>  inp_feat(365), I3 =>  inp_feat(360), I4 =>  inp_feat(436), I5 =>  inp_feat(71), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_52_S_0_L_1_inst : LUT8 generic map(INIT => "1111110011100100101100111010000000110011010000000010011100000000111101010000000000110001000000000111111100000000001101000000000011001101000001010001111100100000000000010000000100110111000000011010000010000000101100010011000000000000000000000000000000000000") port map( O =>C_52_S_0_L_1_out, I0 =>  inp_feat(6), I1 =>  inp_feat(15), I2 =>  inp_feat(23), I3 =>  inp_feat(183), I4 =>  inp_feat(333), I5 =>  inp_feat(373), I6 =>  inp_feat(143), I7 =>  inp_feat(80)); 
C_52_S_0_L_2_inst : LUT8 generic map(INIT => "1110000011001000111000001110000011100000100000001010000001000000101011111110111010101111100010000011001001111010101011111010101000001000101010001010000000000000101000001100000010100000001000001010000001100110101000001010001010000000001000001000000010000010") port map( O =>C_52_S_0_L_2_out, I0 =>  inp_feat(466), I1 =>  inp_feat(480), I2 =>  inp_feat(87), I3 =>  inp_feat(285), I4 =>  inp_feat(317), I5 =>  inp_feat(203), I6 =>  inp_feat(86), I7 =>  inp_feat(71)); 
C_52_S_0_L_3_inst : LUT8 generic map(INIT => "1111110000011100111111001110110011110010101011111111000011111110000011001100110010101100100011001010101010001010101010101001111111111100010100001000110011001000111100000101011100000000010101010000110010000000000011001101100000000000011101000000000011011111") port map( O =>C_52_S_0_L_3_out, I0 =>  inp_feat(154), I1 =>  inp_feat(297), I2 =>  inp_feat(475), I3 =>  inp_feat(428), I4 =>  inp_feat(362), I5 =>  inp_feat(107), I6 =>  inp_feat(310), I7 =>  inp_feat(151)); 
C_52_S_0_L_4_inst : LUT8 generic map(INIT => "1111111111111111001111101111000011111111110010001010101100000000110000001110101010000000100000000000000000000000110010000000000001010010110000001000001010000000011101110000000000000000000000001100000011000000101000000000000000000000000000000000000000000000") port map( O =>C_52_S_0_L_4_out, I0 =>  inp_feat(373), I1 =>  inp_feat(130), I2 =>  inp_feat(183), I3 =>  inp_feat(145), I4 =>  inp_feat(469), I5 =>  inp_feat(5), I6 =>  inp_feat(74), I7 =>  inp_feat(1)); 
C_52_S_0_L_5_inst : LUT8 generic map(INIT => "1011111110100000111110101000101010111011000000001111101100001010000010010000000011110110000000000100000000000000111100000000000011111100110110001110111111001110110000000000000011111010000010101011111110010000111101100100100011110000100000001111110011000000") port map( O =>C_52_S_0_L_5_out, I0 =>  inp_feat(428), I1 =>  inp_feat(220), I2 =>  inp_feat(331), I3 =>  inp_feat(267), I4 =>  inp_feat(304), I5 =>  inp_feat(79), I6 =>  inp_feat(365), I7 =>  inp_feat(340)); 
C_52_S_0_L_6_inst : LUT8 generic map(INIT => "1011111111011010111011110010001111101111111011100110111110101010001000001010000001111111000000000000100000100000000011111000101010111100110000001100011100000001110010000000110001001111000010111010101010100000011101110000000100001100000000000001111100001010") port map( O =>C_52_S_0_L_6_out, I0 =>  inp_feat(216), I1 =>  inp_feat(212), I2 =>  inp_feat(266), I3 =>  inp_feat(365), I4 =>  inp_feat(101), I5 =>  inp_feat(428), I6 =>  inp_feat(12), I7 =>  inp_feat(103)); 
C_52_S_0_L_7_inst : LUT8 generic map(INIT => "1110110111010101110001001011000111101100111111101100010011000100011001001101111100100100111101111110010011000100100001001100010011001100010000001001110111011001110011001110111001000100100100000100010000000100110001000001000101000000010001000100010011010000") port map( O =>C_52_S_0_L_7_out, I0 =>  inp_feat(318), I1 =>  inp_feat(229), I2 =>  inp_feat(328), I3 =>  inp_feat(420), I4 =>  inp_feat(152), I5 =>  inp_feat(367), I6 =>  inp_feat(373), I7 =>  inp_feat(316)); 
C_52_S_1_L_0_inst : LUT8 generic map(INIT => "1110110110110101111101001111110100000000100100001001000011010000101110010101010111111110000111001000100010000000100000101100000011111000110000000100110010000000000000001000000000000000100000000011100011000000111010101000000000000000110000000000000010000000") port map( O =>C_52_S_1_L_0_out, I0 =>  inp_feat(365), I1 =>  inp_feat(427), I2 =>  inp_feat(504), I3 =>  inp_feat(143), I4 =>  inp_feat(328), I5 =>  inp_feat(267), I6 =>  inp_feat(71), I7 =>  inp_feat(80)); 
C_52_S_1_L_1_inst : LUT8 generic map(INIT => "1111111111111111010100100111111011110100110111101111010001000100100100011000111100000000001010111100000000000000000000000000000011010001101110000000000110010001101101110011001011110101111100110001000000000000000000000000000000010001000000000000000000000000") port map( O =>C_52_S_1_L_1_out, I0 =>  inp_feat(494), I1 =>  inp_feat(86), I2 =>  inp_feat(365), I3 =>  inp_feat(340), I4 =>  inp_feat(373), I5 =>  inp_feat(151), I6 =>  inp_feat(60), I7 =>  inp_feat(216)); 
C_52_S_1_L_2_inst : LUT8 generic map(INIT => "1110111011000000111010100010001011100110101000000111101100100010110011000000000010100000000000000000000000000000101110110010001001101011101000101111110111100000101011111010101011111111011001010000000000000000000001010000000000000000000000001011110000000000") port map( O =>C_52_S_1_L_2_out, I0 =>  inp_feat(216), I1 =>  inp_feat(232), I2 =>  inp_feat(87), I3 =>  inp_feat(439), I4 =>  inp_feat(107), I5 =>  inp_feat(100), I6 =>  inp_feat(296), I7 =>  inp_feat(31)); 
C_52_S_1_L_3_inst : LUT8 generic map(INIT => "0010101100000011001100111010111110011000000100001100111111011111101000001000100010100000000000001000100000000000000000000000000011111110101100001111111100000000000000000000000000000000000000001000000000000000101000000000000000000000000000000000000000000000") port map( O =>C_52_S_1_L_3_out, I0 =>  inp_feat(263), I1 =>  inp_feat(317), I2 =>  inp_feat(106), I3 =>  inp_feat(90), I4 =>  inp_feat(101), I5 =>  inp_feat(12), I6 =>  inp_feat(470), I7 =>  inp_feat(378)); 
C_52_S_1_L_4_inst : LUT8 generic map(INIT => "1101101111101101110111011111111111010100000111011100000001001100110111001110110000000100110011000100010011010000000001000000010010001000000011011000001011101110100000000000000000000100000001000000000000000000000000000000000011000000000000000000000000000000") port map( O =>C_52_S_1_L_4_out, I0 =>  inp_feat(362), I1 =>  inp_feat(351), I2 =>  inp_feat(178), I3 =>  inp_feat(367), I4 =>  inp_feat(164), I5 =>  inp_feat(105), I6 =>  inp_feat(310), I7 =>  inp_feat(294)); 
C_52_S_1_L_5_inst : LUT8 generic map(INIT => "1111010111111101101000001000100011111110100000000000000000000000111000001100000010100000100000001111000010000000110000000000000011000000110100000000000001000000110001011000000000000000000000000010000011000000010000001000000011000000110000001100000000000000") port map( O =>C_52_S_1_L_5_out, I0 =>  inp_feat(263), I1 =>  inp_feat(87), I2 =>  inp_feat(54), I3 =>  inp_feat(56), I4 =>  inp_feat(158), I5 =>  inp_feat(220), I6 =>  inp_feat(6), I7 =>  inp_feat(277)); 
C_52_S_1_L_6_inst : LUT8 generic map(INIT => "1101111011011000111111000010110011001100100000000000110000000000110010001000000000001100100001001000110010001000000011000000010011011100010000000111100000000000100001001000000000000000000000001000110000000000000011001000000010001100000000000000000000000000") port map( O =>C_52_S_1_L_6_out, I0 =>  inp_feat(477), I1 =>  inp_feat(296), I2 =>  inp_feat(139), I3 =>  inp_feat(80), I4 =>  inp_feat(5), I5 =>  inp_feat(504), I6 =>  inp_feat(6), I7 =>  inp_feat(310)); 
C_52_S_1_L_7_inst : LUT8 generic map(INIT => "0010101100000000111001000100000011110111100000001111000011101011000000010010000011000000000000001011001000000000111101101110001111100000100000001100110000000000110100011000000011010100110000001000000010000000000000001000000011000000101000001111000010100000") port map( O =>C_52_S_1_L_7_out, I0 =>  inp_feat(267), I1 =>  inp_feat(396), I2 =>  inp_feat(439), I3 =>  inp_feat(365), I4 =>  inp_feat(340), I5 =>  inp_feat(0), I6 =>  inp_feat(87), I7 =>  inp_feat(262)); 
C_52_S_2_L_0_inst : LUT8 generic map(INIT => "1111110001001111111011000010000011100000001000000010100000100000110010100000000010000000000000001100000000000000000000000000000011101100100011100000100010001000000000000000000000101000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_52_S_2_L_0_out, I0 =>  inp_feat(303), I1 =>  inp_feat(80), I2 =>  inp_feat(475), I3 =>  inp_feat(183), I4 =>  inp_feat(101), I5 =>  inp_feat(12), I6 =>  inp_feat(345), I7 =>  inp_feat(216)); 
C_52_S_2_L_1_inst : LUT8 generic map(INIT => "1111110011110100111101111000000011100100000010001111000000000000111111000010010011111101001100000010000000000000010100000000000011000000000000000100100000000000000000001000000010001100000000001100000010001000111111000000100010001000100010001000000000000000") port map( O =>C_52_S_2_L_1_out, I0 =>  inp_feat(317), I1 =>  inp_feat(49), I2 =>  inp_feat(87), I3 =>  inp_feat(201), I4 =>  inp_feat(200), I5 =>  inp_feat(183), I6 =>  inp_feat(64), I7 =>  inp_feat(285)); 
C_52_S_2_L_2_inst : LUT8 generic map(INIT => "1110101111101110101010110010001011101011011011101010001110100000111011100000000000000000000000001000001010001000100000000000000010101111001010100110101100100000100000101000000011100000000000001100010000000000000000000000000010000000000000001000000000000000") port map( O =>C_52_S_2_L_2_out, I0 =>  inp_feat(480), I1 =>  inp_feat(169), I2 =>  inp_feat(221), I3 =>  inp_feat(80), I4 =>  inp_feat(316), I5 =>  inp_feat(42), I6 =>  inp_feat(132), I7 =>  inp_feat(53)); 
C_52_S_2_L_3_inst : LUT8 generic map(INIT => "0000100111101000001010001010100010000010001000000000000010001000110010001110000010100000101000001000000000000000000000000000000011111011111000001000100010101000011110100000000000000000000000001010000010100000000000001010000000000000000000000000000000000000") port map( O =>C_52_S_2_L_3_out, I0 =>  inp_feat(74), I1 =>  inp_feat(63), I2 =>  inp_feat(255), I3 =>  inp_feat(262), I4 =>  inp_feat(296), I5 =>  inp_feat(281), I6 =>  inp_feat(492), I7 =>  inp_feat(151)); 
C_52_S_2_L_4_inst : LUT8 generic map(INIT => "1110000011100000111110101000100011001000101000001110000010111000111001100000000011111000001000001111100010100000111000001010000011111111111100001011100011111000000010000000000000000000111100001111111011100100101110101111000100001000000000000000000000000000") port map( O =>C_52_S_2_L_4_out, I0 =>  inp_feat(103), I1 =>  inp_feat(392), I2 =>  inp_feat(87), I3 =>  inp_feat(33), I4 =>  inp_feat(56), I5 =>  inp_feat(73), I6 =>  inp_feat(203), I7 =>  inp_feat(101)); 
C_52_S_2_L_5_inst : LUT8 generic map(INIT => "1111111110101010000010101010000001101010111000001000000010000000110111111010001011001010000000000010000010000010000000000000000011100010111010101010101010100010000000101000000010000010000000000111101000000010101000100000000000000000000000000000000000000000") port map( O =>C_52_S_2_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(107), I2 =>  inp_feat(297), I3 =>  inp_feat(310), I4 =>  inp_feat(201), I5 =>  inp_feat(477), I6 =>  inp_feat(351), I7 =>  inp_feat(158)); 
C_52_S_2_L_6_inst : LUT8 generic map(INIT => "1111101111111000101101111110111111010101111101001110011011111011101011000000000000000000000000001010110000000000000000000000000011101110101110001000000010100000001010101111110000000000110100000000101100000000000000000000000000000001000000000000000000000000") port map( O =>C_52_S_2_L_6_out, I0 =>  inp_feat(451), I1 =>  inp_feat(251), I2 =>  inp_feat(105), I3 =>  inp_feat(239), I4 =>  inp_feat(310), I5 =>  inp_feat(71), I6 =>  inp_feat(146), I7 =>  inp_feat(331)); 
C_52_S_2_L_7_inst : LUT8 generic map(INIT => "1011101011101010011010001110111011101000101000001110100010000010001000001000101011100000111110100011100010111000110011001000001011101000101010101000110000101010111110000001101011111100101011101110100011100010111010000111101011101010101010001100111000001000") port map( O =>C_52_S_2_L_7_out, I0 =>  inp_feat(87), I1 =>  inp_feat(103), I2 =>  inp_feat(282), I3 =>  inp_feat(186), I4 =>  inp_feat(329), I5 =>  inp_feat(285), I6 =>  inp_feat(203), I7 =>  inp_feat(64)); 
C_52_S_3_L_0_inst : LUT8 generic map(INIT => "1010001011101000111000001111000010101001111110000000000011110000001010000000100011100000000000001000100010001000000000001010000010100000000000001010000010000000101000001010101000000000101000001010100010001000101000001000000010001000100010001000000010000000") port map( O =>C_52_S_3_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(296), I2 =>  inp_feat(267), I3 =>  inp_feat(46), I4 =>  inp_feat(157), I5 =>  inp_feat(99), I6 =>  inp_feat(452), I7 =>  inp_feat(492)); 
C_52_S_3_L_1_inst : LUT8 generic map(INIT => "1111110011111100110100000101000011001100001000001001010100010001111111110101000011110000011100001111001110100000100101010011001000100010110000000000000000000000111000111010000000000000000000000011111010000000100000000000000011101011010100001000000100000000") port map( O =>C_52_S_3_L_1_out, I0 =>  inp_feat(186), I1 =>  inp_feat(282), I2 =>  inp_feat(387), I3 =>  inp_feat(158), I4 =>  inp_feat(33), I5 =>  inp_feat(56), I6 =>  inp_feat(200), I7 =>  inp_feat(71)); 
C_52_S_3_L_2_inst : LUT8 generic map(INIT => "1111101010001010101010001010101011111110100001001010101010000000100010111000110010001000100000001000111110001010100010001000100010110010000000001001100010101010111110110000000010101010000000000000000000000000000000000000000010100010000000000000000000000000") port map( O =>C_52_S_3_L_2_out, I0 =>  inp_feat(183), I1 =>  inp_feat(307), I2 =>  inp_feat(323), I3 =>  inp_feat(139), I4 =>  inp_feat(218), I5 =>  inp_feat(200), I6 =>  inp_feat(49), I7 =>  inp_feat(285)); 
C_52_S_3_L_3_inst : LUT8 generic map(INIT => "1111001110100011101100011011110010100010000100001010111000011010100000001000000010100000000100001000000010000000000000000001000011111111111110110011000011010011000000000001000000000000000100111000100011011000000000000011000100000000000000000000000000010000") port map( O =>C_52_S_3_L_3_out, I0 =>  inp_feat(105), I1 =>  inp_feat(301), I2 =>  inp_feat(373), I3 =>  inp_feat(323), I4 =>  inp_feat(9), I5 =>  inp_feat(111), I6 =>  inp_feat(205), I7 =>  inp_feat(130)); 
C_52_S_3_L_4_inst : LUT8 generic map(INIT => "0011110011010000111101000010000011100000111000001101001011000101111010101110101011101000000011100100100010000000111111111110111111101000101000000000000000000000110000001100000000000000000000001100100011001000000010001000100000000000000000000000000000000000") port map( O =>C_52_S_3_L_4_out, I0 =>  inp_feat(272), I1 =>  inp_feat(203), I2 =>  inp_feat(21), I3 =>  inp_feat(103), I4 =>  inp_feat(186), I5 =>  inp_feat(101), I6 =>  inp_feat(130), I7 =>  inp_feat(151)); 
C_52_S_3_L_5_inst : LUT8 generic map(INIT => "1111111111000100111111110100001011100000011011111100001001101010110000001110001001100000001000101100000011100010111000101110001011000011010000101000001100000010010000111110001101000010010000101100001111100000010000110010001011010011111000101100001110000000") port map( O =>C_52_S_3_L_5_out, I0 =>  inp_feat(15), I1 =>  inp_feat(92), I2 =>  inp_feat(316), I3 =>  inp_feat(365), I4 =>  inp_feat(331), I5 =>  inp_feat(340), I6 =>  inp_feat(327), I7 =>  inp_feat(1)); 
C_52_S_3_L_6_inst : LUT8 generic map(INIT => "1100000110000000101110111011101001010101000000011111101110110111101000101000000000100010000000001000000000000000000000000000000011010101110000001111001100101010111100011000100011010001111100101100000001000000010000000100000000010000000000000100000000000000") port map( O =>C_52_S_3_L_6_out, I0 =>  inp_feat(367), I1 =>  inp_feat(301), I2 =>  inp_feat(428), I3 =>  inp_feat(414), I4 =>  inp_feat(340), I5 =>  inp_feat(53), I6 =>  inp_feat(42), I7 =>  inp_feat(29)); 
C_52_S_3_L_7_inst : LUT8 generic map(INIT => "1111111110001101111111111010111010110000000000001010000010001001011111010000010110111001000011110001000100000001100100010000000011111111100001011111111111101011100000001100000010110100011100000101010100000101111110011011100000000000000000001011000110000000") port map( O =>C_52_S_3_L_7_out, I0 =>  inp_feat(272), I1 =>  inp_feat(263), I2 =>  inp_feat(33), I3 =>  inp_feat(387), I4 =>  inp_feat(48), I5 =>  inp_feat(87), I6 =>  inp_feat(428), I7 =>  inp_feat(216)); 
C_52_S_4_L_0_inst : LUT8 generic map(INIT => "1001101001011110100011001000010011011101010001011110010100000100111011000000110010001100000000001001000000000000000000000000000011100000000000001000100000000000101010000000000010100000000000001111110000000000100011000000000001000000000000000000000000000000") port map( O =>C_52_S_4_L_0_out, I0 =>  inp_feat(301), I1 =>  inp_feat(373), I2 =>  inp_feat(9), I3 =>  inp_feat(111), I4 =>  inp_feat(205), I5 =>  inp_feat(130), I6 =>  inp_feat(262), I7 =>  inp_feat(151)); 
C_52_S_4_L_1_inst : LUT8 generic map(INIT => "1111110001000100111111000100110011111100100000000101000011000000111101100000000011010111111000000000000000000000000000000000000001101101000011001111010110001101110101010000010001010101010101000111111100000000111011011000100100000000000000000100010100000100") port map( O =>C_52_S_4_L_1_out, I0 =>  inp_feat(383), I1 =>  inp_feat(316), I2 =>  inp_feat(259), I3 =>  inp_feat(80), I4 =>  inp_feat(362), I5 =>  inp_feat(116), I6 =>  inp_feat(152), I7 =>  inp_feat(5)); 
C_52_S_4_L_2_inst : LUT8 generic map(INIT => "1011000010101000111101111001110011110010111101111010001111101010101010101000000000000010011000001010000010100000001000101000001011101010110000000000000000000000111000000000000000100000000000001010001011000000000000000000000000000000000000001010001000000000") port map( O =>C_52_S_4_L_2_out, I0 =>  inp_feat(81), I1 =>  inp_feat(307), I2 =>  inp_feat(87), I3 =>  inp_feat(218), I4 =>  inp_feat(386), I5 =>  inp_feat(64), I6 =>  inp_feat(262), I7 =>  inp_feat(151)); 
C_52_S_4_L_3_inst : LUT8 generic map(INIT => "1101110111111000111110011111110010001000100010000000000010001000110011001100000011001000110011001000000000000000000000000000000001000100000000000010000000001100010000001100100010000000000010001111100011001000000000001100010010000000010010001100000011001000") port map( O =>C_52_S_4_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(439), I2 =>  inp_feat(297), I3 =>  inp_feat(433), I4 =>  inp_feat(120), I5 =>  inp_feat(238), I6 =>  inp_feat(179), I7 =>  inp_feat(351)); 
C_52_S_4_L_4_inst : LUT8 generic map(INIT => "0110111010101000110111101000000000101000100000001010100010101000101010001010100010111000101110000000000000000000101100001010000010000000000000001111111100000000000000000000000011001010000000000000000010000000110111001000000000000000000000001100100000000000") port map( O =>C_52_S_4_L_4_out, I0 =>  inp_feat(428), I1 =>  inp_feat(222), I2 =>  inp_feat(316), I3 =>  inp_feat(95), I4 =>  inp_feat(221), I5 =>  inp_feat(54), I6 =>  inp_feat(327), I7 =>  inp_feat(1)); 
C_52_S_4_L_5_inst : LUT8 generic map(INIT => "1101101011100101110001011111110111010100000000001111011111001100111101011000010010100010100010000010010000000000000100000000000011111111111011101111111111111111000000000000001000100010001000111010010010100000001100110010001100000000000000000010000000000010") port map( O =>C_52_S_4_L_5_out, I0 =>  inp_feat(317), I1 =>  inp_feat(323), I2 =>  inp_feat(263), I3 =>  inp_feat(384), I4 =>  inp_feat(9), I5 =>  inp_feat(111), I6 =>  inp_feat(205), I7 =>  inp_feat(130)); 
C_52_S_4_L_6_inst : LUT8 generic map(INIT => "0101010111110100111101001111110011011100111111001111110011111110101100000000000010010000100000000011000000110010001100000011000001100100110101000110110001010000101110001111100100100000001100010000000000000000000100000000000010111000101110000011000000110000") port map( O =>C_52_S_4_L_6_out, I0 =>  inp_feat(317), I1 =>  inp_feat(33), I2 =>  inp_feat(87), I3 =>  inp_feat(473), I4 =>  inp_feat(340), I5 =>  inp_feat(101), I6 =>  inp_feat(12), I7 =>  inp_feat(90)); 
C_52_S_4_L_7_inst : LUT8 generic map(INIT => "1111011110001000101110111010100010110101001100001000000001000000101110110000100000001000000010001011100100001000000010000000100011111010100010000100000001001000011000001100000001000000100000000000110000000000100010001000100010110000000000000000000000001000") port map( O =>C_52_S_4_L_7_out, I0 =>  inp_feat(483), I1 =>  inp_feat(221), I2 =>  inp_feat(494), I3 =>  inp_feat(255), I4 =>  inp_feat(477), I5 =>  inp_feat(351), I6 =>  inp_feat(179), I7 =>  inp_feat(87)); 
C_53_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_1_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_2_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_3_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_53_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000001010000000010000000100010001000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000100000000000000010001000") port map( O =>C_53_S_4_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(10), I2 =>  inp_feat(75), I3 =>  inp_feat(293), I4 =>  inp_feat(260), I5 =>  inp_feat(213), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_54_S_0_L_0_inst : LUT8 generic map(INIT => "1111111111111111110011111011110111000000100000000000000000000000111100001111001100000001111000110000000010000000000000000000000010101100000010010000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_54_S_0_L_0_out, I0 =>  inp_feat(201), I1 =>  inp_feat(229), I2 =>  inp_feat(302), I3 =>  inp_feat(336), I4 =>  inp_feat(333), I5 =>  inp_feat(366), I6 =>  inp_feat(217), I7 =>  inp_feat(111)); 
C_54_S_0_L_1_inst : LUT8 generic map(INIT => "0101010001001000110111110100000001001101010010001101111101000000010011111101000011011111110100000100111111110000101011011101000011111000100010001000000000000000100010001000100000000000000000001100000000000000110000000000000000000000000000000000000000000000") port map( O =>C_54_S_0_L_1_out, I0 =>  inp_feat(492), I1 =>  inp_feat(466), I2 =>  inp_feat(377), I3 =>  inp_feat(254), I4 =>  inp_feat(493), I5 =>  inp_feat(166), I6 =>  inp_feat(143), I7 =>  inp_feat(305)); 
C_54_S_0_L_2_inst : LUT8 generic map(INIT => "1111111000110110110000001111010000000000001100101100000011110010110011101111000010101010101001100000000011111101000000001000000011100000100101001100000000010000000000000000001011000000100000001010000010110011000000001011001000000000100100100000000000110000") port map( O =>C_54_S_0_L_2_out, I0 =>  inp_feat(80), I1 =>  inp_feat(383), I2 =>  inp_feat(210), I3 =>  inp_feat(71), I4 =>  inp_feat(266), I5 =>  inp_feat(267), I6 =>  inp_feat(151), I7 =>  inp_feat(216)); 
C_54_S_0_L_3_inst : LUT8 generic map(INIT => "1110111111000000100000000000000001001101110000000001000000000000111110001010000010111000000010000010110011110000110111000000000010000010100000000010000000000000000000000000000000000000000000000011000000110010001100000000000000000000011000000000000000000000") port map( O =>C_54_S_0_L_3_out, I0 =>  inp_feat(229), I1 =>  inp_feat(178), I2 =>  inp_feat(62), I3 =>  inp_feat(90), I4 =>  inp_feat(297), I5 =>  inp_feat(74), I6 =>  inp_feat(221), I7 =>  inp_feat(368)); 
C_54_S_0_L_4_inst : LUT8 generic map(INIT => "1010001011111000001000001110000011001000111110001000001011010001000000001100000000000000101000001100000011000000000000000000000011111000101100001000000010000000100000001010000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_54_S_0_L_4_out, I0 =>  inp_feat(365), I1 =>  inp_feat(238), I2 =>  inp_feat(183), I3 =>  inp_feat(288), I4 =>  inp_feat(135), I5 =>  inp_feat(396), I6 =>  inp_feat(60), I7 =>  inp_feat(305)); 
C_54_S_0_L_5_inst : LUT8 generic map(INIT => "1101011111101000111101111110000011111111110001001111111111100100011000001000000001000100001000000011000011000000000000001010000001100000100000001110000110000000111101101000000011110100101100101010000010000000000000001111001010100000111000000000000011100000") port map( O =>C_54_S_0_L_5_out, I0 =>  inp_feat(285), I1 =>  inp_feat(323), I2 =>  inp_feat(87), I3 =>  inp_feat(33), I4 =>  inp_feat(64), I5 =>  inp_feat(340), I6 =>  inp_feat(12), I7 =>  inp_feat(54)); 
C_54_S_0_L_6_inst : LUT8 generic map(INIT => "1111110111101100111111010101100011001100110010000000000000001000111001000010000011110000000000000000000000000000000000000000000001100100111001010111000011011100110011010100010001010001110111011010000100000000000000000000000000000000000000000000000000000000") port map( O =>C_54_S_0_L_6_out, I0 =>  inp_feat(15), I1 =>  inp_feat(428), I2 =>  inp_feat(201), I3 =>  inp_feat(422), I4 =>  inp_feat(57), I5 =>  inp_feat(294), I6 =>  inp_feat(214), I7 =>  inp_feat(105)); 
C_54_S_0_L_7_inst : LUT8 generic map(INIT => "1011001111011110010110000101000011111000110110001100000010000000111111111100010111011100000001011111010110000101000100000000000010010000100000000100000000100001100000001100100000000000110000001101010110000101010100000101000010010101100001000100000000000000") port map( O =>C_54_S_0_L_7_out, I0 =>  inp_feat(364), I1 =>  inp_feat(351), I2 =>  inp_feat(477), I3 =>  inp_feat(210), I4 =>  inp_feat(310), I5 =>  inp_feat(448), I6 =>  inp_feat(151), I7 =>  inp_feat(373)); 
C_54_S_1_L_0_inst : LUT8 generic map(INIT => "0100010111011101110010001100101010001100010011001100000001001100100011110000110110000100100001010000110110001101101010001000101011110000100010001100000010000000100000000000000010000000000000000000000000000000000000001010101000000000000000001010000010101010") port map( O =>C_54_S_1_L_0_out, I0 =>  inp_feat(396), I1 =>  inp_feat(439), I2 =>  inp_feat(298), I3 =>  inp_feat(328), I4 =>  inp_feat(288), I5 =>  inp_feat(493), I6 =>  inp_feat(143), I7 =>  inp_feat(305)); 
C_54_S_1_L_1_inst : LUT8 generic map(INIT => "1110100011101000001000000000000010100000101000101010000000000000111000000000000010000000000000001010000000000000100000000000000011001000000000000100110011000000000000000000000011000110101000101100000000000000000000000000000011100000000000001111100011100000") port map( O =>C_54_S_1_L_1_out, I0 =>  inp_feat(480), I1 =>  inp_feat(183), I2 =>  inp_feat(54), I3 =>  inp_feat(452), I4 =>  inp_feat(441), I5 =>  inp_feat(381), I6 =>  inp_feat(79), I7 =>  inp_feat(4)); 
C_54_S_1_L_2_inst : LUT8 generic map(INIT => "1111111111001111110111000000101111111110110010000100110000000001111010000000000000000000000000001000110000000000000011000000000011111111011110101111110000010100100111111000110000000001000000001111000010100000101000001000000010000000100000000000000000000000") port map( O =>C_54_S_1_L_2_out, I0 =>  inp_feat(103), I1 =>  inp_feat(267), I2 =>  inp_feat(278), I3 =>  inp_feat(11), I4 =>  inp_feat(183), I5 =>  inp_feat(285), I6 =>  inp_feat(151), I7 =>  inp_feat(149)); 
C_54_S_1_L_3_inst : LUT8 generic map(INIT => "1111101110101000111110111010000011101000100000001000100000000000001110010010100000001000001000001111100000010000011100000011000000011010101010010110111111101110000000000000000000000000000000000010000000000000101010010000110011110000000000001101000000010000") port map( O =>C_54_S_1_L_3_out, I0 =>  inp_feat(87), I1 =>  inp_feat(479), I2 =>  inp_feat(329), I3 =>  inp_feat(483), I4 =>  inp_feat(303), I5 =>  inp_feat(151), I6 =>  inp_feat(71), I7 =>  inp_feat(11)); 
C_54_S_1_L_4_inst : LUT8 generic map(INIT => "1110110111101100110110101111101010001000000011001100100000000000111100000000000011111111111010101111000000000000110000000000000001101111100011001000100000000000101011110110101010001000000010000110010100100000000000000000000000010111000001010000000000000000") port map( O =>C_54_S_1_L_4_out, I0 =>  inp_feat(323), I1 =>  inp_feat(408), I2 =>  inp_feat(15), I3 =>  inp_feat(428), I4 =>  inp_feat(381), I5 =>  inp_feat(57), I6 =>  inp_feat(79), I7 =>  inp_feat(310)); 
C_54_S_1_L_5_inst : LUT8 generic map(INIT => "1010100011000000100010000000100010101000101010000000100000000000101010101000000010101010000000001010100000000000101010100000000001000100010111001001000011000000110010001111110010100100111000001000001011000000100010001000000000000000110100001110000011110000") port map( O =>C_54_S_1_L_5_out, I0 =>  inp_feat(428), I1 =>  inp_feat(466), I2 =>  inp_feat(198), I3 =>  inp_feat(328), I4 =>  inp_feat(422), I5 =>  inp_feat(57), I6 =>  inp_feat(294), I7 =>  inp_feat(161)); 
C_54_S_1_L_6_inst : LUT8 generic map(INIT => "1110110011001100111010001110000000001100000000000010001010000000111011001010000010101000101000001001000000000000101000001010000011001100010011001010001010100000000001000000000010000010000000000101110110000000111111111111000011011100100000001101101110000000") port map( O =>C_54_S_1_L_6_out, I0 =>  inp_feat(234), I1 =>  inp_feat(373), I2 =>  inp_feat(79), I3 =>  inp_feat(138), I4 =>  inp_feat(340), I5 =>  inp_feat(480), I6 =>  inp_feat(221), I7 =>  inp_feat(105)); 
C_54_S_1_L_7_inst : LUT8 generic map(INIT => "0100101011111010001010110010000111111010000110000010000000000000101010101000101010101111001001111110001000000000001110010000000011101000110010100100000000001010110110000111100001000000000000001000100000000000100011010000111111101100110010001111111100001000") port map( O =>C_54_S_1_L_7_out, I0 =>  inp_feat(322), I1 =>  inp_feat(317), I2 =>  inp_feat(56), I3 =>  inp_feat(218), I4 =>  inp_feat(33), I5 =>  inp_feat(108), I6 =>  inp_feat(106), I7 =>  inp_feat(130)); 
C_54_S_2_L_0_inst : LUT8 generic map(INIT => "1110111000101000111110101110001011101010010000001111101111111111100010101000000010001010100010100000111001000000000010100000001011110000101000001011100010101000111100001110000011111011101100000000000000000000000010100000000011001010000000000000001000000010") port map( O =>C_54_S_2_L_0_out, I0 =>  inp_feat(87), I1 =>  inp_feat(282), I2 =>  inp_feat(33), I3 =>  inp_feat(365), I4 =>  inp_feat(340), I5 =>  inp_feat(64), I6 =>  inp_feat(12), I7 =>  inp_feat(216)); 
C_54_S_2_L_1_inst : LUT8 generic map(INIT => "1111001010101000100000001000000011111110001010101010001100000000111110011111100011000000010000001101110111001000110101010000000010001000001000001011001000001000111100101010000010111000010000001110010111110000101111110111000111001101000000011111110100000000") port map( O =>C_54_S_2_L_1_out, I0 =>  inp_feat(87), I1 =>  inp_feat(362), I2 =>  inp_feat(297), I3 =>  inp_feat(210), I4 =>  inp_feat(267), I5 =>  inp_feat(340), I6 =>  inp_feat(151), I7 =>  inp_feat(504)); 
C_54_S_2_L_2_inst : LUT8 generic map(INIT => "1011111111111011001011111111100101110001011111000011001111000011101111110111111100001011101111000100000000111011000000110000000110111000111110000000100000000000100010000000000000000000000000001110110010001000000010000000000010001000100010000000000000000000") port map( O =>C_54_S_2_L_2_out, I0 =>  inp_feat(115), I1 =>  inp_feat(340), I2 =>  inp_feat(475), I3 =>  inp_feat(29), I4 =>  inp_feat(310), I5 =>  inp_feat(105), I6 =>  inp_feat(316), I7 =>  inp_feat(305)); 
C_54_S_2_L_3_inst : LUT8 generic map(INIT => "1010111000000000111011100010001000001100000000001111110100000000111100001110010011100000111011111100010011101000110100000110101011100000101000101010000010101010000000000000000010100000100000001000000001000000100000001000101100000000000000000000000010100000") port map( O =>C_54_S_2_L_3_out, I0 =>  inp_feat(297), I1 =>  inp_feat(5), I2 =>  inp_feat(387), I3 =>  inp_feat(153), I4 =>  inp_feat(222), I5 =>  inp_feat(373), I6 =>  inp_feat(105), I7 =>  inp_feat(90)); 
C_54_S_2_L_4_inst : LUT8 generic map(INIT => "1011110110111000111101110011100010011000001100100011001100100000100000000010101000100000001000000000000000100000000000000000001010110001101111111110000001110000101000001010001000000000000000000000000010101000001000000000000000000000100000000000000000000000") port map( O =>C_54_S_2_L_4_out, I0 =>  inp_feat(183), I1 =>  inp_feat(383), I2 =>  inp_feat(80), I3 =>  inp_feat(188), I4 =>  inp_feat(216), I5 =>  inp_feat(238), I6 =>  inp_feat(60), I7 =>  inp_feat(296)); 
C_54_S_2_L_5_inst : LUT8 generic map(INIT => "1101110000001100010001001100110011001110110111000111011100011111110111111100010110111011000000111011111110110011101111110011000100001000010000001000100010001100000001011101110100010000000011100101011111001000101010100000001100001110110011111010001000001011") port map( O =>C_54_S_2_L_5_out, I0 =>  inp_feat(52), I1 =>  inp_feat(141), I2 =>  inp_feat(221), I3 =>  inp_feat(316), I4 =>  inp_feat(328), I5 =>  inp_feat(247), I6 =>  inp_feat(261), I7 =>  inp_feat(74)); 
C_54_S_2_L_6_inst : LUT8 generic map(INIT => "0111011100001100011011111110010000111100000110000011110000111000001010000010000000001010001010000000000000100000001010100010101010101100111010001010111000100000101011000000000010101010000000001010100010101000001010100010100000101000000000000010101000000000") port map( O =>C_54_S_2_L_6_out, I0 =>  inp_feat(238), I1 =>  inp_feat(475), I2 =>  inp_feat(178), I3 =>  inp_feat(80), I4 =>  inp_feat(509), I5 =>  inp_feat(271), I6 =>  inp_feat(267), I7 =>  inp_feat(151)); 
C_54_S_2_L_7_inst : LUT8 generic map(INIT => "1101111111110011010010000101111101110110111111110101110010010101110010001100100000000000000000000100000011000000010000000000000000100000101010000000000001000101001011101010001000000000000000001000100010001000000000000000000000000000100000000000000000000000") port map( O =>C_54_S_2_L_7_out, I0 =>  inp_feat(151), I1 =>  inp_feat(298), I2 =>  inp_feat(100), I3 =>  inp_feat(288), I4 =>  inp_feat(135), I5 =>  inp_feat(396), I6 =>  inp_feat(22), I7 =>  inp_feat(60)); 
C_54_S_3_L_0_inst : LUT8 generic map(INIT => "1110110111110010110001011110000011010100110100000101000110000000000010000000000000000001000000001000000000000000000000000000000011101010001000100010001000100000101010100010001000001010001000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_54_S_3_L_0_out, I0 =>  inp_feat(142), I1 =>  inp_feat(413), I2 =>  inp_feat(396), I3 =>  inp_feat(206), I4 =>  inp_feat(105), I5 =>  inp_feat(316), I6 =>  inp_feat(267), I7 =>  inp_feat(305)); 
C_54_S_3_L_1_inst : LUT8 generic map(INIT => "0111011100101000110001001000111010001010100000001010101010100011111011110011010000001111100011111000000000100000101010000001000011100000101000100100000000000000101010100000000010001000000000001110000000000000000000000000000000000000001000000000000000000000") port map( O =>C_54_S_3_L_1_out, I0 =>  inp_feat(23), I1 =>  inp_feat(203), I2 =>  inp_feat(323), I3 =>  inp_feat(71), I4 =>  inp_feat(377), I5 =>  inp_feat(54), I6 =>  inp_feat(285), I7 =>  inp_feat(305)); 
C_54_S_3_L_2_inst : LUT8 generic map(INIT => "1011111011111111011100010111101101110100101000100101000100010001110010001100000000000000100000001000100010000000100000001000000000000000111100100000001011110001000000000100001000000000010100110000000011000000000000000000000000000000110000000000000000000000") port map( O =>C_54_S_3_L_2_out, I0 =>  inp_feat(228), I1 =>  inp_feat(119), I2 =>  inp_feat(120), I3 =>  inp_feat(221), I4 =>  inp_feat(483), I5 =>  inp_feat(331), I6 =>  inp_feat(64), I7 =>  inp_feat(1)); 
C_54_S_3_L_3_inst : LUT8 generic map(INIT => "0110100000001000011000011010000001101000101010001110000110100000000000000000100000000000000000001010000010101010000000000000000011110100000000001011001100100000111010001010100011111111001000000000000000000000000000100010001000000000000010000000001100000010") port map( O =>C_54_S_3_L_3_out, I0 =>  inp_feat(74), I1 =>  inp_feat(30), I2 =>  inp_feat(492), I3 =>  inp_feat(294), I4 =>  inp_feat(178), I5 =>  inp_feat(340), I6 =>  inp_feat(306), I7 =>  inp_feat(247)); 
C_54_S_3_L_4_inst : LUT8 generic map(INIT => "1100100010101010110000001010101011111110101111111100111100100110100100001111101011000000101000101111001011101110110101111111011101000000000000001100010001000000011001100010001001000100101000001000000000000000110000000000000000010000000000001001110011110111") port map( O =>C_54_S_3_L_4_out, I0 =>  inp_feat(161), I1 =>  inp_feat(385), I2 =>  inp_feat(83), I3 =>  inp_feat(82), I4 =>  inp_feat(475), I5 =>  inp_feat(187), I6 =>  inp_feat(316), I7 =>  inp_feat(310)); 
C_54_S_3_L_5_inst : LUT8 generic map(INIT => "0001010111011111101000000000000001100000000000001000000000000000110001000000000000000000000000000000000000000000000000000000000011111110011100010000000000000000110001100000000000000000000000001111111000000001000000000000000000111110000000000000000000000000") port map( O =>C_54_S_3_L_5_out, I0 =>  inp_feat(109), I1 =>  inp_feat(128), I2 =>  inp_feat(480), I3 =>  inp_feat(220), I4 =>  inp_feat(22), I5 =>  inp_feat(306), I6 =>  inp_feat(91), I7 =>  inp_feat(247)); 
C_54_S_3_L_6_inst : LUT8 generic map(INIT => "0110111111111111100111101110111001001100110011010000111011001111101010001000100010100000100000000010000110001000100011101010101011111110100000000110000010000000100000000000000000000000000000001010000000000000000000001000000010001100100010101010101010101010") port map( O =>C_54_S_3_L_6_out, I0 =>  inp_feat(87), I1 =>  inp_feat(365), I2 =>  inp_feat(473), I3 =>  inp_feat(317), I4 =>  inp_feat(71), I5 =>  inp_feat(181), I6 =>  inp_feat(106), I7 =>  inp_feat(12)); 
C_54_S_3_L_7_inst : LUT8 generic map(INIT => "1010111111101111000111101000110111011111111111110001101111101111101100110010001100100000010000001011010101111110000000010111111110101010100000001000000011000000001000000000000000000000000000001010000000000000000000000100000001110001011101010111000101010101") port map( O =>C_54_S_3_L_7_out, I0 =>  inp_feat(268), I1 =>  inp_feat(212), I2 =>  inp_feat(473), I3 =>  inp_feat(317), I4 =>  inp_feat(71), I5 =>  inp_feat(181), I6 =>  inp_feat(106), I7 =>  inp_feat(12)); 
C_54_S_4_L_0_inst : LUT8 generic map(INIT => "0111001111111001111111101110011010101010000000000000101000000010100000111000000010111110011000100000100000000000000010100000001010100000111100001000001010100010001000000000000000000010000000100000000010000000000000000000001000000000000000000000001000000000") port map( O =>C_54_S_4_L_0_out, I0 =>  inp_feat(80), I1 =>  inp_feat(340), I2 =>  inp_feat(427), I3 =>  inp_feat(269), I4 =>  inp_feat(435), I5 =>  inp_feat(242), I6 =>  inp_feat(87), I7 =>  inp_feat(431)); 
C_54_S_4_L_1_inst : LUT8 generic map(INIT => "1111101011110000111100001111000011111110100000101011000011100000111100100000000010110010001000001111101110101010001000100010000011110000100000001010000010000000100010001000000000000000000000001011000000000000101100000010000000111010101000000011001000100000") port map( O =>C_54_S_4_L_1_out, I0 =>  inp_feat(428), I1 =>  inp_feat(222), I2 =>  inp_feat(183), I3 =>  inp_feat(203), I4 =>  inp_feat(139), I5 =>  inp_feat(408), I6 =>  inp_feat(106), I7 =>  inp_feat(277)); 
C_54_S_4_L_2_inst : LUT8 generic map(INIT => "0101111011011111100110000000110111010100110111100100000000001100111111111100111101101100010011001111110011111100010001000000100011001100010001001111000010000000100000001100000000000000000000001000100000001000000000000000000010000000100000000000000000000000") port map( O =>C_54_S_4_L_2_out, I0 =>  inp_feat(195), I1 =>  inp_feat(428), I2 =>  inp_feat(387), I3 =>  inp_feat(322), I4 =>  inp_feat(267), I5 =>  inp_feat(23), I6 =>  inp_feat(130), I7 =>  inp_feat(305)); 
C_54_S_4_L_3_inst : LUT8 generic map(INIT => "1100011010100100111010000000000010111110111000101001100000000000001100001000000011101010000000001110110010001000111110010000000011101100111111001100000001000000110001011111111100000000000000001111110111101000100010000000000011001000110111010000000000000000") port map( O =>C_54_S_4_L_3_out, I0 =>  inp_feat(7), I1 =>  inp_feat(297), I2 =>  inp_feat(267), I3 =>  inp_feat(433), I4 =>  inp_feat(40), I5 =>  inp_feat(176), I6 =>  inp_feat(448), I7 =>  inp_feat(151)); 
C_54_S_4_L_4_inst : LUT8 generic map(INIT => "0010011111101010000010001010101011100010011010101000111011100111011011111000100000001000100010001000000000000000000001000000111111111111111100001000111100000000111111011111000100001111001100101111111110110000000110001000000001110111010101110100111101101011") port map( O =>C_54_S_4_L_4_out, I0 =>  inp_feat(87), I1 =>  inp_feat(232), I2 =>  inp_feat(176), I3 =>  inp_feat(266), I4 =>  inp_feat(267), I5 =>  inp_feat(477), I6 =>  inp_feat(448), I7 =>  inp_feat(151)); 
C_54_S_4_L_5_inst : LUT8 generic map(INIT => "1111011011111110101101100111111111110111110100001001101111010101011100000111101100000000000000000010000000000000000000000000000011001010110010000000100011001000000010100000000000000000000000001100000011111111000000000000000010000000000000000000000000000000") port map( O =>C_54_S_4_L_5_out, I0 =>  inp_feat(304), I1 =>  inp_feat(322), I2 =>  inp_feat(23), I3 =>  inp_feat(0), I4 =>  inp_feat(505), I5 =>  inp_feat(21), I6 =>  inp_feat(306), I7 =>  inp_feat(91)); 
C_54_S_4_L_6_inst : LUT8 generic map(INIT => "1011111010101111001001101010110010110111110101001111101011011100101010000000100000000000000000001001000111010100100011000000010000001000111111100000000011101010010111011101110010001100100011000000111011011101000000000000000011011100110111000000000011001100") port map( O =>C_54_S_4_L_6_out, I0 =>  inp_feat(71), I1 =>  inp_feat(331), I2 =>  inp_feat(6), I3 =>  inp_feat(221), I4 =>  inp_feat(74), I5 =>  inp_feat(210), I6 =>  inp_feat(201), I7 =>  inp_feat(327)); 
C_54_S_4_L_7_inst : LUT8 generic map(INIT => "0001111011100110111010111101011110001000001100100000000000100011101010101000000000111100000000000010000000000000000010000000000011111111001100000010001100010000001111110011101100100010000000111011100000000000001100010000000010101000000001100000000000000010") port map( O =>C_54_S_4_L_7_out, I0 =>  inp_feat(183), I1 =>  inp_feat(80), I2 =>  inp_feat(272), I3 =>  inp_feat(188), I4 =>  inp_feat(5), I5 =>  inp_feat(295), I6 =>  inp_feat(238), I7 =>  inp_feat(0)); 
C_55_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000001010000000000000000000000000000000010000000010110000001100011110101000000000100000000000000010000000000000000000001000000000000010100000000000010000000000000000000100000000010000000011100000101110000000000000000000000000000000000") port map( O =>C_55_S_0_L_0_out, I0 =>  inp_feat(87), I1 =>  inp_feat(109), I2 =>  inp_feat(438), I3 =>  inp_feat(183), I4 =>  inp_feat(267), I5 =>  inp_feat(106), I6 =>  inp_feat(54), I7 =>  inp_feat(111)); 
C_55_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000001000001000000000000000000000000000001000100000010000000000001000100111000100000010100000100010000000000000000111100000000000001011011010100000000000000000000000000000000000000101111000110000001011100000010000000000000000000000000000000000") port map( O =>C_55_S_0_L_1_out, I0 =>  inp_feat(154), I1 =>  inp_feat(267), I2 =>  inp_feat(327), I3 =>  inp_feat(0), I4 =>  inp_feat(387), I5 =>  inp_feat(322), I6 =>  inp_feat(200), I7 =>  inp_feat(71)); 
C_55_S_0_L_2_inst : LUT8 generic map(INIT => "1100000001001100000010000000100001001110000000001000111010001010100011000000000010001000000000001000110100000000100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_0_L_2_out, I0 =>  inp_feat(474), I1 =>  inp_feat(435), I2 =>  inp_feat(428), I3 =>  inp_feat(15), I4 =>  inp_feat(494), I5 =>  inp_feat(87), I6 =>  inp_feat(135), I7 =>  inp_feat(305)); 
C_55_S_0_L_3_inst : LUT8 generic map(INIT => "0000100000000000000010000000000000000000000000000000000000000000000110100000000010001000000000000000000000000000000000000000000010011000000000001000100000000101000000000000000000000000000000000101010000000100100010001100000000000000000000000100010001000000") port map( O =>C_55_S_0_L_3_out, I0 =>  inp_feat(173), I1 =>  inp_feat(266), I2 =>  inp_feat(439), I3 =>  inp_feat(396), I4 =>  inp_feat(310), I5 =>  inp_feat(151), I6 =>  inp_feat(216), I7 =>  inp_feat(437)); 
C_55_S_0_L_4_inst : LUT8 generic map(INIT => "0100100000000000010000000000000010001000010001000001100001000000000000000000000000000000000000000000000000000000000000000000000001011111100011100001111100000000111111111001110100101011000010010000010000000000000000000000000000001101000011000000000000000000") port map( O =>C_55_S_0_L_4_out, I0 =>  inp_feat(272), I1 =>  inp_feat(317), I2 =>  inp_feat(387), I3 =>  inp_feat(9), I4 =>  inp_feat(340), I5 =>  inp_feat(323), I6 =>  inp_feat(12), I7 =>  inp_feat(216)); 
C_55_S_0_L_5_inst : LUT8 generic map(INIT => "1000110001001100000000001000000010010100010001000000000010000000110001000100010100000000000000000101010001000101000000001010000000000000000000000000000000000000000000000000000000000000000000000000000100000101010000000000010000000000000000000000000010100000") port map( O =>C_55_S_0_L_5_out, I0 =>  inp_feat(439), I1 =>  inp_feat(143), I2 =>  inp_feat(428), I3 =>  inp_feat(466), I4 =>  inp_feat(294), I5 =>  inp_feat(385), I6 =>  inp_feat(306), I7 =>  inp_feat(492)); 
C_55_S_0_L_6_inst : LUT8 generic map(INIT => "0000000001000000000001010000010000000000000000000000000000000000000000000100001010001000100011000000000000010000000000001000000011000000100000001000000000000000000000000000000000000000000000001000000011000000010000001100000000000000000000000000000000000000") port map( O =>C_55_S_0_L_6_out, I0 =>  inp_feat(232), I1 =>  inp_feat(151), I2 =>  inp_feat(288), I3 =>  inp_feat(297), I4 =>  inp_feat(80), I5 =>  inp_feat(435), I6 =>  inp_feat(310), I7 =>  inp_feat(316)); 
C_55_S_0_L_7_inst : LUT8 generic map(INIT => "0000010001000000101011100000000000000000000000000000010100000000001000000000000001000000000001000000000000000000000000000000000001000100000000011111000010001101000001001000110110001101000011110000000000000000000000000000000100000000000011000000000000001001") port map( O =>C_55_S_0_L_7_out, I0 =>  inp_feat(90), I1 =>  inp_feat(340), I2 =>  inp_feat(54), I3 =>  inp_feat(15), I4 =>  inp_feat(285), I5 =>  inp_feat(33), I6 =>  inp_feat(473), I7 =>  inp_feat(1)); 
C_55_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000100000000001000000000000000000000000000100001010000000000000000000000000000000000000000010000000000000001010000000000001100000001000000110100000000000011000000000000001111111110101000110010100000000000000000000000001100000000000000") port map( O =>C_55_S_1_L_0_out, I0 =>  inp_feat(310), I1 =>  inp_feat(340), I2 =>  inp_feat(347), I3 =>  inp_feat(20), I4 =>  inp_feat(183), I5 =>  inp_feat(60), I6 =>  inp_feat(160), I7 =>  inp_feat(71)); 
C_55_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000110010101100001111000000000000000100000000000000110000101000000100000000010000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_1_L_1_out, I0 =>  inp_feat(471), I1 =>  inp_feat(224), I2 =>  inp_feat(492), I3 =>  inp_feat(466), I4 =>  inp_feat(316), I5 =>  inp_feat(143), I6 =>  inp_feat(277), I7 =>  inp_feat(305)); 
C_55_S_1_L_2_inst : LUT8 generic map(INIT => "0001000101011000000000000010100000000000000000000000000000001000010100001101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000") port map( O =>C_55_S_1_L_2_out, I0 =>  inp_feat(213), I1 =>  inp_feat(360), I2 =>  inp_feat(218), I3 =>  inp_feat(436), I4 =>  inp_feat(157), I5 =>  inp_feat(73), I6 =>  inp_feat(45), I7 =>  inp_feat(305)); 
C_55_S_1_L_3_inst : LUT8 generic map(INIT => "1001001100001011010000000100001111010001000000110000000000000000000100000101111100000000010101010111100011101111010100000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_1_L_3_out, I0 =>  inp_feat(11), I1 =>  inp_feat(323), I2 =>  inp_feat(33), I3 =>  inp_feat(54), I4 =>  inp_feat(329), I5 =>  inp_feat(87), I6 =>  inp_feat(285), I7 =>  inp_feat(305)); 
C_55_S_1_L_4_inst : LUT8 generic map(INIT => "0001110000000000000001000000000001000100000000000000100000000000010001000000000010000000000000000000000100000000000000000000000010001000000000001011000000000000000011000000000011001100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_1_L_4_out, I0 =>  inp_feat(428), I1 =>  inp_feat(15), I2 =>  inp_feat(466), I3 =>  inp_feat(22), I4 =>  inp_feat(381), I5 =>  inp_feat(332), I6 =>  inp_feat(473), I7 =>  inp_feat(1)); 
C_55_S_1_L_5_inst : LUT8 generic map(INIT => "0010011000011011001011110010001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001100101110000011100110011000000000000000000000001000100000000000000000100000000000000000000000000000000000000000000000000") port map( O =>C_55_S_1_L_5_out, I0 =>  inp_feat(388), I1 =>  inp_feat(87), I2 =>  inp_feat(183), I3 =>  inp_feat(365), I4 =>  inp_feat(281), I5 =>  inp_feat(214), I6 =>  inp_feat(464), I7 =>  inp_feat(238)); 
C_55_S_1_L_6_inst : LUT8 generic map(INIT => "0011101110000000111011010100110100100000000000000010100010101000100000110000000000001100000001001100000000000000000010000010110000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_1_L_6_out, I0 =>  inp_feat(473), I1 =>  inp_feat(183), I2 =>  inp_feat(56), I3 =>  inp_feat(317), I4 =>  inp_feat(370), I5 =>  inp_feat(428), I6 =>  inp_feat(340), I7 =>  inp_feat(12)); 
C_55_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000101000000000000010010000000000001010100000000000000000000000000000000000000000001001000000000000000000000000000010100000000000000111000010010000011100110100000011101000010000100000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_55_S_1_L_7_out, I0 =>  inp_feat(107), I1 =>  inp_feat(494), I2 =>  inp_feat(151), I3 =>  inp_feat(435), I4 =>  inp_feat(310), I5 =>  inp_feat(216), I6 =>  inp_feat(266), I7 =>  inp_feat(373)); 
C_55_S_2_L_0_inst : LUT8 generic map(INIT => "1110001001110011000000000100000100100010111101000000000000000000000000000001000100000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000") port map( O =>C_55_S_2_L_0_out, I0 =>  inp_feat(306), I1 =>  inp_feat(27), I2 =>  inp_feat(61), I3 =>  inp_feat(224), I4 =>  inp_feat(492), I5 =>  inp_feat(471), I6 =>  inp_feat(143), I7 =>  inp_feat(305)); 
C_55_S_2_L_1_inst : LUT8 generic map(INIT => "0000001000001010000010000000100000001010100000000000001000100010101010001000101000000000000010000000000010101010000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_2_L_1_out, I0 =>  inp_feat(40), I1 =>  inp_feat(74), I2 =>  inp_feat(483), I3 =>  inp_feat(87), I4 =>  inp_feat(298), I5 =>  inp_feat(80), I6 =>  inp_feat(431), I7 =>  inp_feat(305)); 
C_55_S_2_L_2_inst : LUT8 generic map(INIT => "0001000000000000001000000000000000000000000000001001000000000000100000000000000010000000000000000000000000000000101100001001000110000000010100000001000000000000010000000000000001110000000000001111010000000000001000000000000100010000000000001111101011111011") port map( O =>C_55_S_2_L_2_out, I0 =>  inp_feat(428), I1 =>  inp_feat(285), I2 =>  inp_feat(473), I3 =>  inp_feat(317), I4 =>  inp_feat(1), I5 =>  inp_feat(33), I6 =>  inp_feat(105), I7 =>  inp_feat(408)); 
C_55_S_2_L_3_inst : LUT8 generic map(INIT => "0000010010000100000000000111110100000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000001100011101001100010110010101000000001001010000000100000001010000000000000100000000000000010100000000000000000000000000000000") port map( O =>C_55_S_2_L_3_out, I0 =>  inp_feat(54), I1 =>  inp_feat(64), I2 =>  inp_feat(71), I3 =>  inp_feat(387), I4 =>  inp_feat(285), I5 =>  inp_feat(340), I6 =>  inp_feat(12), I7 =>  inp_feat(281)); 
C_55_S_2_L_4_inst : LUT8 generic map(INIT => "1010010011100000100010000000000010000000000000001100000110000000101000111000000000001010000000001000000000000000000011010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_2_L_4_out, I0 =>  inp_feat(130), I1 =>  inp_feat(107), I2 =>  inp_feat(6), I3 =>  inp_feat(317), I4 =>  inp_feat(15), I5 =>  inp_feat(138), I6 =>  inp_feat(23), I7 =>  inp_feat(305)); 
C_55_S_2_L_5_inst : LUT8 generic map(INIT => "0001011111000000100000101100000000000000000000000000000000000000111000110100000001110100110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010101000000110000000100000000000000000000000000000101010000") port map( O =>C_55_S_2_L_5_out, I0 =>  inp_feat(480), I1 =>  inp_feat(336), I2 =>  inp_feat(172), I3 =>  inp_feat(466), I4 =>  inp_feat(428), I5 =>  inp_feat(435), I6 =>  inp_feat(310), I7 =>  inp_feat(52)); 
C_55_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000010000000100000001000000000011100101000000000101000100000000010001000110000001000100000001000101010100000000000001000000000010000000000000000000010000000000110001000000001000000000000100000100000001000000000000000000001001000100000000000") port map( O =>C_55_S_2_L_6_out, I0 =>  inp_feat(15), I1 =>  inp_feat(353), I2 =>  inp_feat(344), I3 =>  inp_feat(222), I4 =>  inp_feat(387), I5 =>  inp_feat(183), I6 =>  inp_feat(11), I7 =>  inp_feat(221)); 
C_55_S_2_L_7_inst : LUT8 generic map(INIT => "0000000010001100000000000000000011001000010011000000000000000000110000000100000000000000000001001100000001000100000000000101000000000000000000000000000000000000010000000000000000000000000000000000000100100000000000000000000011010001010101000000000000000100") port map( O =>C_55_S_2_L_7_out, I0 =>  inp_feat(267), I1 =>  inp_feat(151), I2 =>  inp_feat(340), I3 =>  inp_feat(297), I4 =>  inp_feat(435), I5 =>  inp_feat(504), I6 =>  inp_feat(87), I7 =>  inp_feat(288)); 
C_55_S_3_L_0_inst : LUT8 generic map(INIT => "0010000101000000010000000000000010000000000000001100000000000000110000000100000011000000000000001001000000000000110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_55_S_3_L_0_out, I0 =>  inp_feat(306), I1 =>  inp_feat(294), I2 =>  inp_feat(258), I3 =>  inp_feat(227), I4 =>  inp_feat(54), I5 =>  inp_feat(183), I6 =>  inp_feat(90), I7 =>  inp_feat(305)); 
C_55_S_3_L_1_inst : LUT8 generic map(INIT => "1100011100011100000000000000000000100110111000000101001000000000000000000000000000000000000000001000000011110100000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_3_L_1_out, I0 =>  inp_feat(380), I1 =>  inp_feat(316), I2 =>  inp_feat(331), I3 =>  inp_feat(221), I4 =>  inp_feat(227), I5 =>  inp_feat(306), I6 =>  inp_feat(414), I7 =>  inp_feat(305)); 
C_55_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000110000100000101000001010101000011000000000101001100000000000000000000000000000000000000000000000100000001000000010111000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_3_L_2_out, I0 =>  inp_feat(317), I1 =>  inp_feat(267), I2 =>  inp_feat(222), I3 =>  inp_feat(297), I4 =>  inp_feat(195), I5 =>  inp_feat(23), I6 =>  inp_feat(322), I7 =>  inp_feat(305)); 
C_55_S_3_L_3_inst : LUT8 generic map(INIT => "0001000100000010000000001000000011001000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000010000110010001001011000001000100110010000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_3_L_3_out, I0 =>  inp_feat(302), I1 =>  inp_feat(371), I2 =>  inp_feat(428), I3 =>  inp_feat(15), I4 =>  inp_feat(81), I5 =>  inp_feat(23), I6 =>  inp_feat(305), I7 =>  inp_feat(11)); 
C_55_S_3_L_4_inst : LUT8 generic map(INIT => "1010000000000000000010000000010010001100000000010001000100000100000000000000010001001100000011000100010001001100111011100100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_3_L_4_out, I0 =>  inp_feat(203), I1 =>  inp_feat(340), I2 =>  inp_feat(33), I3 =>  inp_feat(97), I4 =>  inp_feat(71), I5 =>  inp_feat(323), I6 =>  inp_feat(285), I7 =>  inp_feat(305)); 
C_55_S_3_L_5_inst : LUT8 generic map(INIT => "1110110100000100000000000000000000010000000011000000000000000000011100001101001000100000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010000000000000000000000000000000000000000000000000") port map( O =>C_55_S_3_L_5_out, I0 =>  inp_feat(373), I1 =>  inp_feat(198), I2 =>  inp_feat(347), I3 =>  inp_feat(306), I4 =>  inp_feat(112), I5 =>  inp_feat(328), I6 =>  inp_feat(224), I7 =>  inp_feat(492)); 
C_55_S_3_L_6_inst : LUT8 generic map(INIT => "0101000000010000000100000000000000110000011100010011001000000000000100000000000010010000000000001101000001000000001100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_55_S_3_L_6_out, I0 =>  inp_feat(135), I1 =>  inp_feat(439), I2 =>  inp_feat(435), I3 =>  inp_feat(396), I4 =>  inp_feat(27), I5 =>  inp_feat(297), I6 =>  inp_feat(285), I7 =>  inp_feat(315)); 
C_55_S_3_L_7_inst : LUT8 generic map(INIT => "0011111101100010001000100000100000000000000000000000000000000000000100000111000000000000000100000000000000000000000000000000000001010111110000000010001000000000001001000000000000000000000000000010010000000000000000000100000000000000000000000000010000000000") port map( O =>C_55_S_3_L_7_out, I0 =>  inp_feat(353), I1 =>  inp_feat(480), I2 =>  inp_feat(259), I3 =>  inp_feat(339), I4 =>  inp_feat(109), I5 =>  inp_feat(227), I6 =>  inp_feat(221), I7 =>  inp_feat(161)); 
C_55_S_4_L_0_inst : LUT8 generic map(INIT => "0000000110000010000000000000000001001100001011110000000000000000000000000010000100000000000000001000010000000101000000000000000011110110000001010100000000000000010001000000010000000000000000000000010100000101000000000000000000000100000011000000000000000000") port map( O =>C_55_S_4_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(53), I2 =>  inp_feat(54), I3 =>  inp_feat(387), I4 =>  inp_feat(328), I5 =>  inp_feat(428), I6 =>  inp_feat(102), I7 =>  inp_feat(160)); 
C_55_S_4_L_1_inst : LUT8 generic map(INIT => "1010001110111111101000101100001000100000110100001010000001011001110100000100000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_4_L_1_out, I0 =>  inp_feat(142), I1 =>  inp_feat(373), I2 =>  inp_feat(41), I3 =>  inp_feat(74), I4 =>  inp_feat(327), I5 =>  inp_feat(247), I6 =>  inp_feat(52), I7 =>  inp_feat(305)); 
C_55_S_4_L_2_inst : LUT8 generic map(INIT => "0110001010000001100010100001010101000000000000000000001000000000000100000000000000000011000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_55_S_4_L_2_out, I0 =>  inp_feat(233), I1 =>  inp_feat(216), I2 =>  inp_feat(33), I3 =>  inp_feat(15), I4 =>  inp_feat(54), I5 =>  inp_feat(30), I6 =>  inp_feat(329), I7 =>  inp_feat(305)); 
C_55_S_4_L_3_inst : LUT8 generic map(INIT => "1000000000111100001100001111000001110000101100000000000000010000011010010000010000010000000000001100000011100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000") port map( O =>C_55_S_4_L_3_out, I0 =>  inp_feat(290), I1 =>  inp_feat(198), I2 =>  inp_feat(328), I3 =>  inp_feat(428), I4 =>  inp_feat(52), I5 =>  inp_feat(54), I6 =>  inp_feat(58), I7 =>  inp_feat(305)); 
C_55_S_4_L_4_inst : LUT8 generic map(INIT => "1000010000000000010011000000000010000101001000000000011000001100110000000000000011000011000010000100011100000000110011110000110000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000001000") port map( O =>C_55_S_4_L_4_out, I0 =>  inp_feat(373), I1 =>  inp_feat(210), I2 =>  inp_feat(380), I3 =>  inp_feat(328), I4 =>  inp_feat(420), I5 =>  inp_feat(390), I6 =>  inp_feat(316), I7 =>  inp_feat(91)); 
C_55_S_4_L_5_inst : LUT8 generic map(INIT => "1000101000000000000000000000000010001000000000000000000000000000000010000100110001001100000000000000100000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000100011001000010011000000000010001000000000000000000000000000") port map( O =>C_55_S_4_L_5_out, I0 =>  inp_feat(383), I1 =>  inp_feat(435), I2 =>  inp_feat(310), I3 =>  inp_feat(328), I4 =>  inp_feat(441), I5 =>  inp_feat(452), I6 =>  inp_feat(437), I7 =>  inp_feat(238)); 
C_55_S_4_L_6_inst : LUT8 generic map(INIT => "1010001000000000001000000000000011010011000000000011000000010000001000000000000010100000000000000010100000000000001100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_55_S_4_L_6_out, I0 =>  inp_feat(340), I1 =>  inp_feat(439), I2 =>  inp_feat(396), I3 =>  inp_feat(239), I4 =>  inp_feat(27), I5 =>  inp_feat(297), I6 =>  inp_feat(285), I7 =>  inp_feat(315)); 
C_55_S_4_L_7_inst : LUT8 generic map(INIT => "0000010010000100000001001000010010000101000011000000000010000000000001001100010011000100010001000000000010000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_55_S_4_L_7_out, I0 =>  inp_feat(439), I1 =>  inp_feat(396), I2 =>  inp_feat(436), I3 =>  inp_feat(344), I4 =>  inp_feat(21), I5 =>  inp_feat(390), I6 =>  inp_feat(316), I7 =>  inp_feat(91)); 
C_56_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_0_out, I0 =>  inp_feat(302), I1 =>  inp_feat(57), I2 =>  inp_feat(396), I3 =>  inp_feat(37), I4 =>  inp_feat(242), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_56_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000101000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_56_S_0_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(478), I2 =>  inp_feat(242), I3 =>  inp_feat(190), I4 =>  inp_feat(418), I5 =>  inp_feat(483), I6 =>  inp_feat(329), I7 =>  inp_feat(375)); 
C_56_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000001000001000010000100000000000000000000001000000000000000010010001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_2_out, I0 =>  inp_feat(265), I1 =>  inp_feat(137), I2 =>  inp_feat(478), I3 =>  inp_feat(152), I4 =>  inp_feat(226), I5 =>  inp_feat(483), I6 =>  inp_feat(224), I7 =>  inp_feat(437)); 
C_56_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_3_out, I0 =>  inp_feat(265), I1 =>  inp_feat(139), I2 =>  inp_feat(467), I3 =>  inp_feat(474), I4 =>  inp_feat(249), I5 =>  inp_feat(450), I6 =>  inp_feat(356), I7 =>  inp_feat(171)); 
C_56_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(408), I2 =>  inp_feat(229), I3 =>  inp_feat(478), I4 =>  inp_feat(424), I5 =>  inp_feat(284), I6 =>  inp_feat(157), I7 =>  inp_feat(488)); 
C_56_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000100000000000000010100001101000001010000000000000000000000010000010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_5_out, I0 =>  inp_feat(329), I1 =>  inp_feat(416), I2 =>  inp_feat(473), I3 =>  inp_feat(227), I4 =>  inp_feat(483), I5 =>  inp_feat(272), I6 =>  inp_feat(203), I7 =>  inp_feat(242)); 
C_56_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000010000001000100011000011001000000010001000101000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_6_out, I0 =>  inp_feat(478), I1 =>  inp_feat(321), I2 =>  inp_feat(75), I3 =>  inp_feat(91), I4 =>  inp_feat(152), I5 =>  inp_feat(437), I6 =>  inp_feat(130), I7 =>  inp_feat(436)); 
C_56_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100101110000001100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000010000000011000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_0_L_7_out, I0 =>  inp_feat(469), I1 =>  inp_feat(473), I2 =>  inp_feat(291), I3 =>  inp_feat(236), I4 =>  inp_feat(476), I5 =>  inp_feat(483), I6 =>  inp_feat(190), I7 =>  inp_feat(201)); 
C_56_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_1_L_0_out, I0 =>  inp_feat(302), I1 =>  inp_feat(57), I2 =>  inp_feat(396), I3 =>  inp_feat(37), I4 =>  inp_feat(242), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_56_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000101000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_56_S_1_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(478), I2 =>  inp_feat(242), I3 =>  inp_feat(190), I4 =>  inp_feat(418), I5 =>  inp_feat(483), I6 =>  inp_feat(329), I7 =>  inp_feat(375)); 
C_56_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000001000001000010000100000000000000000000001000000000000000010010001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_1_L_2_out, I0 =>  inp_feat(265), I1 =>  inp_feat(137), I2 =>  inp_feat(478), I3 =>  inp_feat(152), I4 =>  inp_feat(226), I5 =>  inp_feat(483), I6 =>  inp_feat(224), I7 =>  inp_feat(437)); 
C_56_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_1_L_3_out, I0 =>  inp_feat(265), I1 =>  inp_feat(139), I2 =>  inp_feat(467), I3 =>  inp_feat(474), I4 =>  inp_feat(249), I5 =>  inp_feat(450), I6 =>  inp_feat(356), I7 =>  inp_feat(171)); 
C_56_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000001000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000010101000101010001010100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_1_L_4_out, I0 =>  inp_feat(483), I1 =>  inp_feat(229), I2 =>  inp_feat(478), I3 =>  inp_feat(193), I4 =>  inp_feat(290), I5 =>  inp_feat(284), I6 =>  inp_feat(157), I7 =>  inp_feat(488)); 
C_56_S_1_L_5_inst : LUT8 generic map(INIT => "0110000000000000000000000000000011000000000000000000000000000000110000101000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_1_L_5_out, I0 =>  inp_feat(441), I1 =>  inp_feat(317), I2 =>  inp_feat(465), I3 =>  inp_feat(37), I4 =>  inp_feat(293), I5 =>  inp_feat(38), I6 =>  inp_feat(152), I7 =>  inp_feat(190)); 
C_56_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000111000000000000000000000000000000010000000000000000000001000000010100000000000000000000000000000000000000000000000000000100000001000000000000000000000000010000010100000000000000000000010000000101000000000000000000000") port map( O =>C_56_S_1_L_6_out, I0 =>  inp_feat(195), I1 =>  inp_feat(201), I2 =>  inp_feat(322), I3 =>  inp_feat(488), I4 =>  inp_feat(190), I5 =>  inp_feat(380), I6 =>  inp_feat(437), I7 =>  inp_feat(193)); 
C_56_S_1_L_7_inst : LUT8 generic map(INIT => "0000110000000100000000000000000000000000000001000000000000000000000001000000000000000000000000000000000010000000000000000000000001111101101001000000000010000000000000001010010000000000000000000100000000000000000000000000000000000000100000000000000000000000") port map( O =>C_56_S_1_L_7_out, I0 =>  inp_feat(90), I1 =>  inp_feat(229), I2 =>  inp_feat(437), I3 =>  inp_feat(328), I4 =>  inp_feat(436), I5 =>  inp_feat(91), I6 =>  inp_feat(478), I7 =>  inp_feat(152)); 
C_56_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_2_L_0_out, I0 =>  inp_feat(302), I1 =>  inp_feat(57), I2 =>  inp_feat(396), I3 =>  inp_feat(37), I4 =>  inp_feat(242), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_56_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000101000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_56_S_2_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(478), I2 =>  inp_feat(242), I3 =>  inp_feat(190), I4 =>  inp_feat(418), I5 =>  inp_feat(483), I6 =>  inp_feat(329), I7 =>  inp_feat(375)); 
C_56_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000001000000000000000000010001000100010000000000010000000000010001000100000000000100000000000000010001000") port map( O =>C_56_S_2_L_2_out, I0 =>  inp_feat(322), I1 =>  inp_feat(190), I2 =>  inp_feat(494), I3 =>  inp_feat(483), I4 =>  inp_feat(329), I5 =>  inp_feat(318), I6 =>  inp_feat(193), I7 =>  inp_feat(437)); 
C_56_S_2_L_3_inst : LUT8 generic map(INIT => "0000000011001100000000000000110000000000000010000000010011001100000000000000100000000000010011000000000000000000000011000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_2_L_3_out, I0 =>  inp_feat(114), I1 =>  inp_feat(408), I2 =>  inp_feat(442), I3 =>  inp_feat(483), I4 =>  inp_feat(335), I5 =>  inp_feat(362), I6 =>  inp_feat(201), I7 =>  inp_feat(288)); 
C_56_S_2_L_4_inst : LUT8 generic map(INIT => "0000111100100011000000110000001100000000000000100000100000000000000000100000001000000000000000000000000000000000000000000000000000001000000100010000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_2_L_4_out, I0 =>  inp_feat(201), I1 =>  inp_feat(488), I2 =>  inp_feat(476), I3 =>  inp_feat(336), I4 =>  inp_feat(280), I5 =>  inp_feat(489), I6 =>  inp_feat(130), I7 =>  inp_feat(399)); 
C_56_S_2_L_5_inst : LUT8 generic map(INIT => "0011001000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000") port map( O =>C_56_S_2_L_5_out, I0 =>  inp_feat(322), I1 =>  inp_feat(171), I2 =>  inp_feat(195), I3 =>  inp_feat(403), I4 =>  inp_feat(130), I5 =>  inp_feat(489), I6 =>  inp_feat(436), I7 =>  inp_feat(399)); 
C_56_S_2_L_6_inst : LUT8 generic map(INIT => "0010001100000010001000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100010000000000000000000000000000000000000000000100000000000100010000000100000000000000000000000000000000000") port map( O =>C_56_S_2_L_6_out, I0 =>  inp_feat(130), I1 =>  inp_feat(335), I2 =>  inp_feat(308), I3 =>  inp_feat(229), I4 =>  inp_feat(475), I5 =>  inp_feat(190), I6 =>  inp_feat(132), I7 =>  inp_feat(254)); 
C_56_S_2_L_7_inst : LUT8 generic map(INIT => "0001101101010111000000000000000000010000000000000000000000000000001000101010001000000000000000000000000000001000000000000000000011010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_2_L_7_out, I0 =>  inp_feat(441), I1 =>  inp_feat(172), I2 =>  inp_feat(308), I3 =>  inp_feat(475), I4 =>  inp_feat(190), I5 =>  inp_feat(387), I6 =>  inp_feat(254), I7 =>  inp_feat(284)); 
C_56_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_3_L_0_out, I0 =>  inp_feat(302), I1 =>  inp_feat(57), I2 =>  inp_feat(396), I3 =>  inp_feat(37), I4 =>  inp_feat(242), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_56_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000101000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_56_S_3_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(478), I2 =>  inp_feat(242), I3 =>  inp_feat(190), I4 =>  inp_feat(418), I5 =>  inp_feat(483), I6 =>  inp_feat(329), I7 =>  inp_feat(375)); 
C_56_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000001000000000001000000000000000100010000000000000001000100000001000100000000000100000001000000010001000") port map( O =>C_56_S_3_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(242), I2 =>  inp_feat(494), I3 =>  inp_feat(329), I4 =>  inp_feat(488), I5 =>  inp_feat(318), I6 =>  inp_feat(193), I7 =>  inp_feat(437)); 
C_56_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000111010000000000000000000001010001100100000000000000000000000000000000000000000000000000000101000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000") port map( O =>C_56_S_3_L_3_out, I0 =>  inp_feat(7), I1 =>  inp_feat(483), I2 =>  inp_feat(375), I3 =>  inp_feat(301), I4 =>  inp_feat(249), I5 =>  inp_feat(418), I6 =>  inp_feat(405), I7 =>  inp_feat(399)); 
C_56_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000001100000000000000010000000000000101000000000000000000000000000000010000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000") port map( O =>C_56_S_3_L_4_out, I0 =>  inp_feat(488), I1 =>  inp_feat(335), I2 =>  inp_feat(445), I3 =>  inp_feat(157), I4 =>  inp_feat(329), I5 =>  inp_feat(483), I6 =>  inp_feat(221), I7 =>  inp_feat(322)); 
C_56_S_3_L_5_inst : LUT8 generic map(INIT => "1000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_3_L_5_out, I0 =>  inp_feat(157), I1 =>  inp_feat(288), I2 =>  inp_feat(130), I3 =>  inp_feat(137), I4 =>  inp_feat(269), I5 =>  inp_feat(304), I6 =>  inp_feat(242), I7 =>  inp_feat(190)); 
C_56_S_3_L_6_inst : LUT8 generic map(INIT => "0101011100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_3_L_6_out, I0 =>  inp_feat(467), I1 =>  inp_feat(114), I2 =>  inp_feat(172), I3 =>  inp_feat(473), I4 =>  inp_feat(57), I5 =>  inp_feat(242), I6 =>  inp_feat(332), I7 =>  inp_feat(478)); 
C_56_S_3_L_7_inst : LUT8 generic map(INIT => "0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000010000000000000001000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_3_L_7_out, I0 =>  inp_feat(143), I1 =>  inp_feat(476), I2 =>  inp_feat(46), I3 =>  inp_feat(422), I4 =>  inp_feat(473), I5 =>  inp_feat(242), I6 =>  inp_feat(478), I7 =>  inp_feat(488)); 
C_56_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_4_L_0_out, I0 =>  inp_feat(302), I1 =>  inp_feat(57), I2 =>  inp_feat(396), I3 =>  inp_feat(37), I4 =>  inp_feat(242), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_56_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000101000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_56_S_4_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(478), I2 =>  inp_feat(242), I3 =>  inp_feat(190), I4 =>  inp_feat(418), I5 =>  inp_feat(483), I6 =>  inp_feat(329), I7 =>  inp_feat(375)); 
C_56_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100010000000100010001000000000000000000000000000100010000000000000000000000000001000000010000000000000001000000000001000") port map( O =>C_56_S_4_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(242), I2 =>  inp_feat(494), I3 =>  inp_feat(488), I4 =>  inp_feat(442), I5 =>  inp_feat(480), I6 =>  inp_feat(284), I7 =>  inp_feat(437)); 
C_56_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000111010000000000000000000001010001100100000000000000000000000000000000000000000000000000000101000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000") port map( O =>C_56_S_4_L_3_out, I0 =>  inp_feat(7), I1 =>  inp_feat(483), I2 =>  inp_feat(375), I3 =>  inp_feat(301), I4 =>  inp_feat(338), I5 =>  inp_feat(418), I6 =>  inp_feat(405), I7 =>  inp_feat(399)); 
C_56_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000100000000000000010000000100000001000011110000000000000000000000000100100000000001000000000000000100000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000") port map( O =>C_56_S_4_L_4_out, I0 =>  inp_feat(437), I1 =>  inp_feat(184), I2 =>  inp_feat(291), I3 =>  inp_feat(222), I4 =>  inp_feat(483), I5 =>  inp_feat(108), I6 =>  inp_feat(221), I7 =>  inp_feat(322)); 
C_56_S_4_L_5_inst : LUT8 generic map(INIT => "1100101010000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_4_L_5_out, I0 =>  inp_feat(271), I1 =>  inp_feat(465), I2 =>  inp_feat(317), I3 =>  inp_feat(378), I4 =>  inp_feat(130), I5 =>  inp_feat(242), I6 =>  inp_feat(304), I7 =>  inp_feat(190)); 
C_56_S_4_L_6_inst : LUT8 generic map(INIT => "0100000000001001000000000000000001011100000000000000000100010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_4_L_6_out, I0 =>  inp_feat(222), I1 =>  inp_feat(170), I2 =>  inp_feat(416), I3 =>  inp_feat(317), I4 =>  inp_feat(479), I5 =>  inp_feat(152), I6 =>  inp_feat(190), I7 =>  inp_feat(408)); 
C_56_S_4_L_7_inst : LUT8 generic map(INIT => "0001000000000000000000000000000000000000000000000000000000000000011101010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_56_S_4_L_7_out, I0 =>  inp_feat(467), I1 =>  inp_feat(416), I2 =>  inp_feat(478), I3 =>  inp_feat(494), I4 =>  inp_feat(398), I5 =>  inp_feat(190), I6 =>  inp_feat(171), I7 =>  inp_feat(37)); 
C_57_S_0_L_0_inst : LUT8 generic map(INIT => "1110111011101010101000001100000011001100100000001010000010000000100011001100000010000000110000001100100011000000110000001000000000000010000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000110000001000000010000000") port map( O =>C_57_S_0_L_0_out, I0 =>  inp_feat(115), I1 =>  inp_feat(375), I2 =>  inp_feat(305), I3 =>  inp_feat(324), I4 =>  inp_feat(60), I5 =>  inp_feat(387), I6 =>  inp_feat(264), I7 =>  inp_feat(488)); 
C_57_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_0_L_2_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_0_L_3_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_0_L_4_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_0_L_5_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_0_L_6_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_0_L_7_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_0_inst : LUT8 generic map(INIT => "1110111011101010101000001100000011001100100000001010000010000000100011001100000010000000110000001100100011000000110000001000000000000010000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000110000001000000010000000") port map( O =>C_57_S_1_L_0_out, I0 =>  inp_feat(115), I1 =>  inp_feat(375), I2 =>  inp_feat(305), I3 =>  inp_feat(324), I4 =>  inp_feat(60), I5 =>  inp_feat(387), I6 =>  inp_feat(264), I7 =>  inp_feat(488)); 
C_57_S_1_L_1_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_2_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_3_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_4_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_5_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_6_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_1_L_7_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_1_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_0_inst : LUT8 generic map(INIT => "1110111011101010101000001100000011001100100000001010000010000000100011001100000010000000110000001100100011000000110000001000000000000010000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000110000001000000010000000") port map( O =>C_57_S_2_L_0_out, I0 =>  inp_feat(115), I1 =>  inp_feat(375), I2 =>  inp_feat(305), I3 =>  inp_feat(324), I4 =>  inp_feat(60), I5 =>  inp_feat(387), I6 =>  inp_feat(264), I7 =>  inp_feat(488)); 
C_57_S_2_L_1_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_2_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_3_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_4_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_5_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_6_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_2_L_7_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_2_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_0_inst : LUT8 generic map(INIT => "1110111011101010101000001100000011001100100000001010000010000000100011001100000010000000110000001100100011000000110000001000000000000010000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000110000001000000010000000") port map( O =>C_57_S_3_L_0_out, I0 =>  inp_feat(115), I1 =>  inp_feat(375), I2 =>  inp_feat(305), I3 =>  inp_feat(324), I4 =>  inp_feat(60), I5 =>  inp_feat(387), I6 =>  inp_feat(264), I7 =>  inp_feat(488)); 
C_57_S_3_L_1_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_2_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_3_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_4_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_5_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_6_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_3_L_7_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_3_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_0_inst : LUT8 generic map(INIT => "1110111011101010101000001100000011001100100000001010000010000000100011001100000010000000110000001100100011000000110000001000000000000010000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000110000001000000010000000") port map( O =>C_57_S_4_L_0_out, I0 =>  inp_feat(115), I1 =>  inp_feat(375), I2 =>  inp_feat(305), I3 =>  inp_feat(324), I4 =>  inp_feat(60), I5 =>  inp_feat(387), I6 =>  inp_feat(264), I7 =>  inp_feat(488)); 
C_57_S_4_L_1_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_2_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_3_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_4_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_5_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_6_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_57_S_4_L_7_inst : LUT8 generic map(INIT => "1111111111111111111110111001010111110010111000001000000000000000000000010000100100010001000100010000000000000000000000000000000011111000111011011011000010110011000100000000000000000000000000000011000000000001000100010000000100000000000000000000000000000000") port map( O =>C_57_S_4_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(222), I3 =>  inp_feat(190), I4 =>  inp_feat(60), I5 =>  inp_feat(476), I6 =>  inp_feat(488), I7 =>  inp_feat(483)); 
C_58_S_0_L_0_inst : LUT8 generic map(INIT => "1111110011000000111101001100000011101100110101001111110011000000101111001010001100110000000000000001100011011000000000000000000000000000010000000101010001000000010011000100010011010100010101000000000000000000000000000000000000000000000000000000000000010000") port map( O =>C_58_S_0_L_0_out, I0 =>  inp_feat(171), I1 =>  inp_feat(226), I2 =>  inp_feat(256), I3 =>  inp_feat(152), I4 =>  inp_feat(322), I5 =>  inp_feat(190), I6 =>  inp_feat(204), I7 =>  inp_feat(488)); 
C_58_S_0_L_1_inst : LUT8 generic map(INIT => "1111111111111110111111111100110011101110110011000000000000000000101011100000101011010110110010000010111001000000000000000100000011101110111011100000110100000100111000100000000000000000000000000000001000000010000000000000000000000000000000000000000000000000") port map( O =>C_58_S_0_L_1_out, I0 =>  inp_feat(473), I1 =>  inp_feat(352), I2 =>  inp_feat(307), I3 =>  inp_feat(237), I4 =>  inp_feat(329), I5 =>  inp_feat(459), I6 =>  inp_feat(115), I7 =>  inp_feat(483)); 
C_58_S_0_L_2_inst : LUT8 generic map(INIT => "1111111110100000111111011100000001001000010001000100010001000000110010001000000000000000000000001100100010001000000000000000000011000000100000000100000011000000010010000000000001000000000000001100100010000000000000000000000011001000000000000000000000000000") port map( O =>C_58_S_0_L_2_out, I0 =>  inp_feat(372), I1 =>  inp_feat(226), I2 =>  inp_feat(152), I3 =>  inp_feat(114), I4 =>  inp_feat(444), I5 =>  inp_feat(416), I6 =>  inp_feat(209), I7 =>  inp_feat(437)); 
C_58_S_0_L_3_inst : LUT8 generic map(INIT => "1010111110101010110010110000000011000001100010010100001000000000111011111010101111110111000000001111111111111111110001010000000011100111110000001110001000000000101000001000000000100010000000001111010100000000100000000000000001010000100000000000000000000000") port map( O =>C_58_S_0_L_3_out, I0 =>  inp_feat(283), I1 =>  inp_feat(290), I2 =>  inp_feat(87), I3 =>  inp_feat(256), I4 =>  inp_feat(475), I5 =>  inp_feat(130), I6 =>  inp_feat(190), I7 =>  inp_feat(288)); 
C_58_S_0_L_4_inst : LUT8 generic map(INIT => "1110100011101110101011011111111111001000101011001010000011111111000000000010100010100100101111011000000010101000000000001111100100000000000000000010000000100000111011000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_0_L_4_out, I0 =>  inp_feat(128), I1 =>  inp_feat(444), I2 =>  inp_feat(242), I3 =>  inp_feat(478), I4 =>  inp_feat(473), I5 =>  inp_feat(130), I6 =>  inp_feat(483), I7 =>  inp_feat(335)); 
C_58_S_0_L_5_inst : LUT8 generic map(INIT => "1110111111111000111011001011100001001100000000001111110010110000110011111000000010101000101010000000100000100000100010001001100011100000101000001000000000000000000000000000000010100000000000000010000010000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_0_L_5_out, I0 =>  inp_feat(475), I1 =>  inp_feat(128), I2 =>  inp_feat(444), I3 =>  inp_feat(437), I4 =>  inp_feat(474), I5 =>  inp_feat(459), I6 =>  inp_feat(483), I7 =>  inp_feat(75)); 
C_58_S_0_L_6_inst : LUT8 generic map(INIT => "1111101101001010110000100100001001110000000000000000000000000000111111110000001011110111000000101111000100000000001000000000000011111000111110101100000011010000111110100101000000000000000000000111111100000000010111010000000011110101000100000000010100000000") port map( O =>C_58_S_0_L_6_out, I0 =>  inp_feat(422), I1 =>  inp_feat(130), I2 =>  inp_feat(387), I3 =>  inp_feat(437), I4 =>  inp_feat(128), I5 =>  inp_feat(152), I6 =>  inp_feat(274), I7 =>  inp_feat(436)); 
C_58_S_0_L_7_inst : LUT8 generic map(INIT => "1111101111111000111111101111000110100010000000000010000000000000111000110000000011100011000000001111001000000000100000000000000010101000101100001010100011100000000000000000000000000000000000001011001110110000000000000000000011110111011101100000000000000000") port map( O =>C_58_S_0_L_7_out, I0 =>  inp_feat(398), I1 =>  inp_feat(478), I2 =>  inp_feat(475), I3 =>  inp_feat(483), I4 =>  inp_feat(437), I5 =>  inp_feat(329), I6 =>  inp_feat(509), I7 =>  inp_feat(217)); 
C_58_S_1_L_0_inst : LUT8 generic map(INIT => "1111110011000000111101001100000011101100110101001111110011000000101111001010001100110000000000000001100011011000000000000000000000000000010000000101010001000000010011000100010011010100010101000000000000000000000000000000000000000000000000000000000000010000") port map( O =>C_58_S_1_L_0_out, I0 =>  inp_feat(171), I1 =>  inp_feat(226), I2 =>  inp_feat(256), I3 =>  inp_feat(152), I4 =>  inp_feat(322), I5 =>  inp_feat(190), I6 =>  inp_feat(204), I7 =>  inp_feat(488)); 
C_58_S_1_L_1_inst : LUT8 generic map(INIT => "0011000011111100111000001110000011000000010000001100000011000000111100001011000011000000100000000000000000000000100000000000000011110111111111110000000010100000100000000000000011001100000000000011000000110000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_1_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(242), I2 =>  inp_feat(488), I3 =>  inp_feat(61), I4 =>  inp_feat(474), I5 =>  inp_feat(508), I6 =>  inp_feat(288), I7 =>  inp_feat(387)); 
C_58_S_1_L_2_inst : LUT8 generic map(INIT => "1111111111001110110011111101101100001100000000001000111000000000110011000100000011001100110000000000100000000000100011000000000010001000100010000000000010000000000000000000000000001000000000000000000010000000000010001000000000001000000000001100100000000000") port map( O =>C_58_S_1_L_2_out, I0 =>  inp_feat(483), I1 =>  inp_feat(488), I2 =>  inp_feat(478), I3 =>  inp_feat(91), I4 =>  inp_feat(100), I5 =>  inp_feat(255), I6 =>  inp_feat(437), I7 =>  inp_feat(476)); 
C_58_S_1_L_3_inst : LUT8 generic map(INIT => "1111110011111111100000001110110010000000011011001000000010100000000010001101111110001000000010000000100010000100000010001000100010101010101011110000000000000000000000000000000000000000000000000000110011001100000000000000100000001000010011000000000000001000") port map( O =>C_58_S_1_L_3_out, I0 =>  inp_feat(444), I1 =>  inp_feat(152), I2 =>  inp_feat(408), I3 =>  inp_feat(478), I4 =>  inp_feat(325), I5 =>  inp_feat(115), I6 =>  inp_feat(128), I7 =>  inp_feat(439)); 
C_58_S_1_L_4_inst : LUT8 generic map(INIT => "1111111111111100111011101010111010000000111000000000000000000000000111011010101011101111100011100010000000000000000000000000000011011100101000001000110000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_1_L_4_out, I0 =>  inp_feat(419), I1 =>  inp_feat(256), I2 =>  inp_feat(87), I3 =>  inp_feat(130), I4 =>  inp_feat(398), I5 =>  inp_feat(335), I6 =>  inp_feat(483), I7 =>  inp_feat(226)); 
C_58_S_1_L_5_inst : LUT8 generic map(INIT => "1111001011110010111100000011001011110011001110110101010111111111111100011011000011000000000000001111001101110010000000000000000010100000000000000000000000000000101101111010000100000100000000101110000011000000000000000000000011100010110000010000000000000000") port map( O =>C_58_S_1_L_5_out, I0 =>  inp_feat(307), I1 =>  inp_feat(190), I2 =>  inp_feat(488), I3 =>  inp_feat(444), I4 =>  inp_feat(128), I5 =>  inp_feat(57), I6 =>  inp_feat(136), I7 =>  inp_feat(226)); 
C_58_S_1_L_6_inst : LUT8 generic map(INIT => "1111110111111010111011101111011111110000110000001100000011110100110010001000000010000000111000001000000010000000000000001100000010101000000000001010000000000000000000000000000000000000000000001100100010000000100000000000000000000000000000001000000010000000") port map( O =>C_58_S_1_L_6_out, I0 =>  inp_feat(475), I1 =>  inp_feat(444), I2 =>  inp_feat(483), I3 =>  inp_feat(143), I4 =>  inp_feat(329), I5 =>  inp_feat(226), I6 =>  inp_feat(288), I7 =>  inp_feat(418)); 
C_58_S_1_L_7_inst : LUT8 generic map(INIT => "1111111010000000111111001111101010001000000000000100010000000000100000000000000011100000010000001000000000000000000000001000000011111111111010101111111010011111100010001000000001000100110011000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_1_L_7_out, I0 =>  inp_feat(130), I1 =>  inp_feat(483), I2 =>  inp_feat(437), I3 =>  inp_feat(256), I4 =>  inp_feat(108), I5 =>  inp_feat(418), I6 =>  inp_feat(226), I7 =>  inp_feat(265)); 
C_58_S_2_L_0_inst : LUT8 generic map(INIT => "1111110011000000111101001100000011101100110101001111110011000000101111001010001100110000000000000001100011011000000000000000000000000000010000000101010001000000010011000100010011010100010101000000000000000000000000000000000000000000000000000000000000010000") port map( O =>C_58_S_2_L_0_out, I0 =>  inp_feat(171), I1 =>  inp_feat(226), I2 =>  inp_feat(256), I3 =>  inp_feat(152), I4 =>  inp_feat(322), I5 =>  inp_feat(190), I6 =>  inp_feat(204), I7 =>  inp_feat(488)); 
C_58_S_2_L_1_inst : LUT8 generic map(INIT => "0101111000100000111110100000000010110000000000001011000000000000111011100000000010100000000000000000000000000000101000000000000011111111001111111000101000000000110000000000000000110000001100000000111100000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_2_L_1_out, I0 =>  inp_feat(256), I1 =>  inp_feat(190), I2 =>  inp_feat(242), I3 =>  inp_feat(488), I4 =>  inp_feat(474), I5 =>  inp_feat(508), I6 =>  inp_feat(288), I7 =>  inp_feat(387)); 
C_58_S_2_L_2_inst : LUT8 generic map(INIT => "1100100000010100111100000100000011110000111100000000000000000000101000001110000010000000111011000000000010000000000000000000000011000000111001001100010001000000000000001111000000000000000000001000000011000100000000001100010000000000110000000000000000000000") port map( O =>C_58_S_2_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(476), I2 =>  inp_feat(488), I3 =>  inp_feat(478), I4 =>  inp_feat(83), I5 =>  inp_feat(156), I6 =>  inp_feat(87), I7 =>  inp_feat(195)); 
C_58_S_2_L_3_inst : LUT8 generic map(INIT => "1101110111011100100011001010100011001101100000000000000000000000110101000000000000000000000000000100000000000000000000000000000011110100111100000000000000000000000001001100000000000000000000001101010001000000000000000000000011001100000000000000000000000000") port map( O =>C_58_S_2_L_3_out, I0 =>  inp_feat(479), I1 =>  inp_feat(488), I2 =>  inp_feat(351), I3 =>  inp_feat(152), I4 =>  inp_feat(375), I5 =>  inp_feat(115), I6 =>  inp_feat(128), I7 =>  inp_feat(32)); 
C_58_S_2_L_4_inst : LUT8 generic map(INIT => "1010101011101010101110100010101011100000111011101010101000101010100010000000101000001010000010100000000000000000000000000000100010000010001000101010001000000010000000000000000000000000000000101010000000000000001000100000000000000000000000000000000000000000") port map( O =>C_58_S_2_L_4_out, I0 =>  inp_feat(488), I1 =>  inp_feat(80), I2 =>  inp_feat(290), I3 =>  inp_feat(87), I4 =>  inp_feat(338), I5 =>  inp_feat(483), I6 =>  inp_feat(179), I7 =>  inp_feat(476)); 
C_58_S_2_L_5_inst : LUT8 generic map(INIT => "1111111111111011110011001000100010100000101010100000000010000000101110101011000110001000100010001010000000100000100000001000100000001110010100110000000010001000000000000000000000000000100000001100100000000000100000001000000000000000000000000000000000000000") port map( O =>C_58_S_2_L_5_out, I0 =>  inp_feat(242), I1 =>  inp_feat(73), I2 =>  inp_feat(130), I3 =>  inp_feat(3), I4 =>  inp_feat(120), I5 =>  inp_feat(476), I6 =>  inp_feat(267), I7 =>  inp_feat(483)); 
C_58_S_2_L_6_inst : LUT8 generic map(INIT => "1111111110111101110111111010100011101111000000001100010010000000110111111000110001001110101010100001111110001000000010100000000011111111101011010000110100000000000000010000000000000000000000000010111100000100000000000000000000001111000000000000000000000000") port map( O =>C_58_S_2_L_6_out, I0 =>  inp_feat(444), I1 =>  inp_feat(130), I2 =>  inp_feat(376), I3 =>  inp_feat(418), I4 =>  inp_feat(459), I5 =>  inp_feat(483), I6 =>  inp_feat(307), I7 =>  inp_feat(329)); 
C_58_S_2_L_7_inst : LUT8 generic map(INIT => "1111110011101000111111101010110011001010000000000000000000000000100010100000000010000000000000001000100000000000000000000000000010100000101010001010000010101000000000000000000000000000000000000000100000000000000000000000000000101000000000000000000000000000") port map( O =>C_58_S_2_L_7_out, I0 =>  inp_feat(459), I1 =>  inp_feat(418), I2 =>  inp_feat(199), I3 =>  inp_feat(238), I4 =>  inp_feat(437), I5 =>  inp_feat(226), I6 =>  inp_feat(152), I7 =>  inp_feat(256)); 
C_58_S_3_L_0_inst : LUT8 generic map(INIT => "1111110011000000111101001100000011101100110101001111110011000000101111001010001100110000000000000001100011011000000000000000000000000000010000000101010001000000010011000100010011010100010101000000000000000000000000000000000000000000000000000000000000010000") port map( O =>C_58_S_3_L_0_out, I0 =>  inp_feat(171), I1 =>  inp_feat(226), I2 =>  inp_feat(256), I3 =>  inp_feat(152), I4 =>  inp_feat(322), I5 =>  inp_feat(190), I6 =>  inp_feat(204), I7 =>  inp_feat(488)); 
C_58_S_3_L_1_inst : LUT8 generic map(INIT => "0101111000100000111110100000000010110000000000001011000000000000111011100000000010100000000000000000000000000000101000000000000011111111001111111000101000000000110000000000000000110000001100000000111100000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_3_L_1_out, I0 =>  inp_feat(256), I1 =>  inp_feat(190), I2 =>  inp_feat(242), I3 =>  inp_feat(488), I4 =>  inp_feat(474), I5 =>  inp_feat(508), I6 =>  inp_feat(288), I7 =>  inp_feat(387)); 
C_58_S_3_L_2_inst : LUT8 generic map(INIT => "1110101111111011111000101100000010101000110001001100100011001000110010001110100011001000111010000100000011000100010010001100010011101010111000001110101010101010000000000100000011101000110000000000000000100000111010101010100000000000000000001000100010000000") port map( O =>C_58_S_3_L_2_out, I0 =>  inp_feat(437), I1 =>  inp_feat(152), I2 =>  inp_feat(475), I3 =>  inp_feat(436), I4 =>  inp_feat(478), I5 =>  inp_feat(272), I6 =>  inp_feat(87), I7 =>  inp_feat(195)); 
C_58_S_3_L_3_inst : LUT8 generic map(INIT => "1111101011111010100010001000100011111010111010101100100000000000001000000000000011001000000000001100000000000000110010100000000000100000101000001000000000000000111100000010000011000000000000001000000000000000100000000000000011000000000000001100000000000000") port map( O =>C_58_S_3_L_3_out, I0 =>  inp_feat(416), I1 =>  inp_feat(29), I2 =>  inp_feat(226), I3 =>  inp_feat(152), I4 =>  inp_feat(216), I5 =>  inp_feat(372), I6 =>  inp_feat(213), I7 =>  inp_feat(483)); 
C_58_S_3_L_4_inst : LUT8 generic map(INIT => "1111100110110111100010100000000010101100000010010000000000000000101110111011101110101010000000000101001000111011000000000000000011111000101000001010100000100000101100000000000010000000000000001101000001000000000000000000000001010000000100000000000000000000") port map( O =>C_58_S_3_L_4_out, I0 =>  inp_feat(444), I1 =>  inp_feat(478), I2 =>  inp_feat(273), I3 =>  inp_feat(509), I4 =>  inp_feat(476), I5 =>  inp_feat(483), I6 =>  inp_feat(61), I7 =>  inp_feat(338)); 
C_58_S_3_L_5_inst : LUT8 generic map(INIT => "1110111011101100100010000000000010101000111010000010000000000000100000001100111000000000000000001010000011001110000000000000000010100000111011000000000000000000001000000000000000000000000000001111101011101110000000000000000011001110111011000000000000000000") port map( O =>C_58_S_3_L_5_out, I0 =>  inp_feat(91), I1 =>  inp_feat(475), I2 =>  inp_feat(329), I3 =>  inp_feat(61), I4 =>  inp_feat(279), I5 =>  inp_feat(444), I6 =>  inp_feat(176), I7 =>  inp_feat(3)); 
C_58_S_3_L_6_inst : LUT8 generic map(INIT => "1110101110001010100010100000100010001000000000001000000000000000111010111010101110101011001010001010101100100010100000100010000010101010101000000000000000000000000000000000000000000000100000001110101100101010100010100000100000000000001000000000000000000000") port map( O =>C_58_S_3_L_6_out, I0 =>  inp_feat(488), I1 =>  inp_feat(142), I2 =>  inp_feat(372), I3 =>  inp_feat(430), I4 =>  inp_feat(504), I5 =>  inp_feat(226), I6 =>  inp_feat(478), I7 =>  inp_feat(256)); 
C_58_S_3_L_7_inst : LUT8 generic map(INIT => "1011110111100100111100100000000011100000100000001110000000000000101011111010110110110011101000001010000000100000101000101000000010110010000000000011001100000000101000001000000000000000000000001010100000100010101110110000100010101010101000001010100000101010") port map( O =>C_58_S_3_L_7_out, I0 =>  inp_feat(383), I1 =>  inp_feat(130), I2 =>  inp_feat(128), I3 =>  inp_feat(483), I4 =>  inp_feat(242), I5 =>  inp_feat(445), I6 =>  inp_feat(379), I7 =>  inp_feat(139)); 
C_58_S_4_L_0_inst : LUT8 generic map(INIT => "1111110011000000111101001100000011101100110101001111110011000000101111001010001100110000000000000001100011011000000000000000000000000000010000000101010001000000010011000100010011010100010101000000000000000000000000000000000000000000000000000000000000010000") port map( O =>C_58_S_4_L_0_out, I0 =>  inp_feat(171), I1 =>  inp_feat(226), I2 =>  inp_feat(256), I3 =>  inp_feat(152), I4 =>  inp_feat(322), I5 =>  inp_feat(190), I6 =>  inp_feat(204), I7 =>  inp_feat(488)); 
C_58_S_4_L_1_inst : LUT8 generic map(INIT => "0101111000100000111110100000000010110000000000001011000000000000111011100000000010100000000000000000000000000000101000000000000011111111001111111000101000000000110000000000000000110000001100000000111100000000000000000000000000000000000000000000000000000000") port map( O =>C_58_S_4_L_1_out, I0 =>  inp_feat(256), I1 =>  inp_feat(190), I2 =>  inp_feat(242), I3 =>  inp_feat(488), I4 =>  inp_feat(474), I5 =>  inp_feat(508), I6 =>  inp_feat(288), I7 =>  inp_feat(387)); 
C_58_S_4_L_2_inst : LUT8 generic map(INIT => "1110101111111011111000101100000010101000110001001100100011001000110010001110100011001000111010000100000011000100010010001100010011101010111000001110101010101010000000000100000011101000110000000000000000100000111010101010100000000000000000001000100010000000") port map( O =>C_58_S_4_L_2_out, I0 =>  inp_feat(437), I1 =>  inp_feat(152), I2 =>  inp_feat(475), I3 =>  inp_feat(436), I4 =>  inp_feat(478), I5 =>  inp_feat(272), I6 =>  inp_feat(87), I7 =>  inp_feat(195)); 
C_58_S_4_L_3_inst : LUT8 generic map(INIT => "1111101011111010100010001000100011111010111010101100100000000000001000000000000011001000000000001100000000000000110010100000000000100000101000001000000000000000111100000010000011000000000000001000000000000000100000000000000011000000000000001100000000000000") port map( O =>C_58_S_4_L_3_out, I0 =>  inp_feat(416), I1 =>  inp_feat(29), I2 =>  inp_feat(226), I3 =>  inp_feat(152), I4 =>  inp_feat(216), I5 =>  inp_feat(372), I6 =>  inp_feat(213), I7 =>  inp_feat(483)); 
C_58_S_4_L_4_inst : LUT8 generic map(INIT => "1001101111001111001000010000101111010001110011000000000000000000101011110000111110101010000010111010011100000000000000000000000011111111010101111010011100000000101001110100010110000000000000001010001100000000000000000000000010000001000000000000000000000000") port map( O =>C_58_S_4_L_4_out, I0 =>  inp_feat(307), I1 =>  inp_feat(298), I2 =>  inp_feat(478), I3 =>  inp_feat(216), I4 =>  inp_feat(476), I5 =>  inp_feat(483), I6 =>  inp_feat(61), I7 =>  inp_feat(338)); 
C_58_S_4_L_5_inst : LUT8 generic map(INIT => "1111111011001100111010001000000000111100100110001111011111100010010000000000000010100000100010000000000100000000101000010000000011110001010101011010000010000000010101010101010101110011111101110111000000000000000000000000000000010101000000010100011100110110") port map( O =>C_58_S_4_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(100), I2 =>  inp_feat(322), I3 =>  inp_feat(29), I4 =>  inp_feat(37), I5 =>  inp_feat(142), I6 =>  inp_feat(128), I7 =>  inp_feat(422)); 
C_58_S_4_L_6_inst : LUT8 generic map(INIT => "1111111111000000111100111000100010100000110010001010000010001000111011111100010011111111101111001010100010000000101110001011111111110000000000001000000011000000100000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_58_S_4_L_6_out, I0 =>  inp_feat(483), I1 =>  inp_feat(94), I2 =>  inp_feat(256), I3 =>  inp_feat(444), I4 =>  inp_feat(171), I5 =>  inp_feat(139), I6 =>  inp_feat(467), I7 =>  inp_feat(375)); 
C_58_S_4_L_7_inst : LUT8 generic map(INIT => "1111111011011000000110000101100011000000111100000000000000110000110010001100100010001000100010000000000000000000000000000000000011111000110110001001000011011000100000000000000000000000100000000110000010000000000000001000000000000000000000000000000000000000") port map( O =>C_58_S_4_L_7_out, I0 =>  inp_feat(87), I1 =>  inp_feat(308), I2 =>  inp_feat(152), I3 =>  inp_feat(270), I4 =>  inp_feat(375), I5 =>  inp_feat(442), I6 =>  inp_feat(173), I7 =>  inp_feat(351)); 
C_59_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000111000001000000000000000010000000100000001000000000000000000000000000000000000000000000000000000010000000100000") port map( O =>C_59_S_0_L_0_out, I0 =>  inp_feat(476), I1 =>  inp_feat(6), I2 =>  inp_feat(431), I3 =>  inp_feat(207), I4 =>  inp_feat(187), I5 =>  inp_feat(79), I6 =>  inp_feat(100), I7 =>  inp_feat(488)); 
C_59_S_0_L_1_inst : LUT8 generic map(INIT => "0101000000000000000000000000000001110000000000000000000000000000101100000000000011110000000000000001000000000000000000000000000000000000000000000000000000000000111100100000000000100010000000000000000000000000000000100000000011111010000000000010101000000000") port map( O =>C_59_S_0_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(475), I2 =>  inp_feat(397), I3 =>  inp_feat(457), I4 =>  inp_feat(66), I5 =>  inp_feat(476), I6 =>  inp_feat(414), I7 =>  inp_feat(375)); 
C_59_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000010000000000000101000000000000000100000100000001010000000000000000000000000000000000000000000000000000010001010101000000000000010000000000000000000000000000000000010000000001000100000100000001000000000000000000010000000000000000000000000101010") port map( O =>C_59_S_0_L_2_out, I0 =>  inp_feat(359), I1 =>  inp_feat(166), I2 =>  inp_feat(176), I3 =>  inp_feat(177), I4 =>  inp_feat(272), I5 =>  inp_feat(437), I6 =>  inp_feat(347), I7 =>  inp_feat(261)); 
C_59_S_0_L_3_inst : LUT8 generic map(INIT => "1000000000001010001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101010101010101110001111001100000000000000100000101010100000000000000000001010000000001000000000000000000000000000000000") port map( O =>C_59_S_0_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(11), I2 =>  inp_feat(500), I3 =>  inp_feat(184), I4 =>  inp_feat(341), I5 =>  inp_feat(224), I6 =>  inp_feat(219), I7 =>  inp_feat(468)); 
C_59_S_0_L_4_inst : LUT8 generic map(INIT => "0101010000001100000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010100000001000000000000000000010011011010101000000000000010000000000000000000000000000000000001000100000010000000000000000000") port map( O =>C_59_S_0_L_4_out, I0 =>  inp_feat(440), I1 =>  inp_feat(100), I2 =>  inp_feat(11), I3 =>  inp_feat(51), I4 =>  inp_feat(224), I5 =>  inp_feat(341), I6 =>  inp_feat(219), I7 =>  inp_feat(292)); 
C_59_S_0_L_5_inst : LUT8 generic map(INIT => "0000000001000100001000000100000000000000010010000110000001100000000100101000001011100100110011000000000000000000111011000110010000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100010000000000000000000100010011000000") port map( O =>C_59_S_0_L_5_out, I0 =>  inp_feat(309), I1 =>  inp_feat(418), I2 =>  inp_feat(473), I3 =>  inp_feat(158), I4 =>  inp_feat(476), I5 =>  inp_feat(177), I6 =>  inp_feat(362), I7 =>  inp_feat(431)); 
C_59_S_0_L_6_inst : LUT8 generic map(INIT => "0101010000001000000000000000000011001110000001010000000000000000001011010000010000000000000000000100111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000001000001011010000000000000000") port map( O =>C_59_S_0_L_6_out, I0 =>  inp_feat(488), I1 =>  inp_feat(23), I2 =>  inp_feat(290), I3 =>  inp_feat(137), I4 =>  inp_feat(277), I5 =>  inp_feat(416), I6 =>  inp_feat(222), I7 =>  inp_feat(61)); 
C_59_S_0_L_7_inst : LUT8 generic map(INIT => "1100001100000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001011100110000000000000000000001010001010100000101000100010000001010100011000000000000000000000000000000000000000000000000") port map( O =>C_59_S_0_L_7_out, I0 =>  inp_feat(51), I1 =>  inp_feat(11), I2 =>  inp_feat(184), I3 =>  inp_feat(411), I4 =>  inp_feat(224), I5 =>  inp_feat(112), I6 =>  inp_feat(22), I7 =>  inp_feat(292)); 
C_59_S_1_L_0_inst : LUT8 generic map(INIT => "0001000000000000110011000001000000000000000000000000000000000000000010100100110111101111010011010000000000000000000000100000000010000010000000000000100000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000000000000") port map( O =>C_59_S_1_L_0_out, I0 =>  inp_feat(222), I1 =>  inp_feat(23), I2 =>  inp_feat(416), I3 =>  inp_feat(478), I4 =>  inp_feat(488), I5 =>  inp_feat(457), I6 =>  inp_feat(239), I7 =>  inp_feat(164)); 
C_59_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000101010000000001000000000000000000000000000000000000000001000000000000000100000000000000000000000000000100010000000000000001010100100000000100000000000000010001000101000001010000000001010101000000000000010000000000000011010000000000000101") port map( O =>C_59_S_1_L_1_out, I0 =>  inp_feat(4), I1 =>  inp_feat(158), I2 =>  inp_feat(177), I3 =>  inp_feat(369), I4 =>  inp_feat(380), I5 =>  inp_feat(459), I6 =>  inp_feat(347), I7 =>  inp_feat(476)); 
C_59_S_1_L_2_inst : LUT8 generic map(INIT => "0010000000000000000000000000000000100000001000100000000000000000101000100000000000000000000000000000000000000000000000000000000001100010100000000000000000000000000000000000000000000000000000001110001000100000010000000000000001000000000000000000000000000000") port map( O =>C_59_S_1_L_2_out, I0 =>  inp_feat(107), I1 =>  inp_feat(418), I2 =>  inp_feat(130), I3 =>  inp_feat(7), I4 =>  inp_feat(471), I5 =>  inp_feat(224), I6 =>  inp_feat(184), I7 =>  inp_feat(441)); 
C_59_S_1_L_3_inst : LUT8 generic map(INIT => "0100000000000000000000000000000001000000001000000000000000010000000000001000000000100000000000100001000000000010011100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000111000000100010") port map( O =>C_59_S_1_L_3_out, I0 =>  inp_feat(440), I1 =>  inp_feat(459), I2 =>  inp_feat(112), I3 =>  inp_feat(51), I4 =>  inp_feat(11), I5 =>  inp_feat(468), I6 =>  inp_feat(341), I7 =>  inp_feat(219)); 
C_59_S_1_L_4_inst : LUT8 generic map(INIT => "0010001000000000111100000010000000101100000000000110110010100000000000000000000000000000000000000000010000000000000000000000000010100100100000000101000001110000001001000000000000110100101000000000000000000000000000000000000000000100000000000000000000000000") port map( O =>C_59_S_1_L_4_out, I0 =>  inp_feat(190), I1 =>  inp_feat(483), I2 =>  inp_feat(497), I3 =>  inp_feat(387), I4 =>  inp_feat(358), I5 =>  inp_feat(475), I6 =>  inp_feat(431), I7 =>  inp_feat(182)); 
C_59_S_1_L_5_inst : LUT8 generic map(INIT => "1100000000000000100110000000000000010000000000000001000000000000000000000000000000000000000000000011010000000000001100110000010000110000000000000000010000000000100111000000000010010001100000000100000010000000000000000000000011010000100000001101000010000000") port map( O =>C_59_S_1_L_5_out, I0 =>  inp_feat(483), I1 =>  inp_feat(53), I2 =>  inp_feat(478), I3 =>  inp_feat(411), I4 =>  inp_feat(6), I5 =>  inp_feat(468), I6 =>  inp_feat(11), I7 =>  inp_feat(459)); 
C_59_S_1_L_6_inst : LUT8 generic map(INIT => "0011000000000000001000000000001000000000000000001010000000000000000000000000000000101000000000001010000010000000101000000000000000000000000000000010000000000000000000000000000000100000000000000000000010000000001000000000010000000000110000001010000000000000") port map( O =>C_59_S_1_L_6_out, I0 =>  inp_feat(100), I1 =>  inp_feat(483), I2 =>  inp_feat(338), I3 =>  inp_feat(474), I4 =>  inp_feat(418), I5 =>  inp_feat(459), I6 =>  inp_feat(441), I7 =>  inp_feat(280)); 
C_59_S_1_L_7_inst : LUT8 generic map(INIT => "0001000001000101010001010100010100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000101010101011100010101000101011000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_1_L_7_out, I0 =>  inp_feat(4), I1 =>  inp_feat(378), I2 =>  inp_feat(436), I3 =>  inp_feat(158), I4 =>  inp_feat(475), I5 =>  inp_feat(270), I6 =>  inp_feat(89), I7 =>  inp_feat(177)); 
C_59_S_2_L_0_inst : LUT8 generic map(INIT => "0000000010100000000010000000000000100011111000000100101100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_2_L_0_out, I0 =>  inp_feat(100), I1 =>  inp_feat(469), I2 =>  inp_feat(107), I3 =>  inp_feat(418), I4 =>  inp_feat(132), I5 =>  inp_feat(139), I6 =>  inp_feat(61), I7 =>  inp_feat(277)); 
C_59_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000010000001100000000000000000000000100000011000000001000000100000000000000010100000000000000000000000000001100000000000000010000000100000001000001100000000000000001000000110000100000000010100000000100000001000000000000000000000000000010000000") port map( O =>C_59_S_2_L_1_out, I0 =>  inp_feat(193), I1 =>  inp_feat(23), I2 =>  inp_feat(377), I3 =>  inp_feat(114), I4 =>  inp_feat(440), I5 =>  inp_feat(449), I6 =>  inp_feat(414), I7 =>  inp_feat(362)); 
C_59_S_2_L_2_inst : LUT8 generic map(INIT => "0001101100100010000000000010001001110011011100110000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_2_L_2_out, I0 =>  inp_feat(56), I1 =>  inp_feat(4), I2 =>  inp_feat(158), I3 =>  inp_feat(475), I4 =>  inp_feat(45), I5 =>  inp_feat(177), I6 =>  inp_feat(457), I7 =>  inp_feat(277)); 
C_59_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000101001101000000000000000000000000000000000000000000001000000011100010010001000000000000000000000000000011010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000") port map( O =>C_59_S_2_L_3_out, I0 =>  inp_feat(11), I1 =>  inp_feat(112), I2 =>  inp_feat(496), I3 =>  inp_feat(280), I4 =>  inp_feat(441), I5 =>  inp_feat(50), I6 =>  inp_feat(184), I7 =>  inp_feat(219)); 
C_59_S_2_L_4_inst : LUT8 generic map(INIT => "0010000000000000000000000000000000000000001000001010000000000000000000000010000000000000000000001100000010110000110011001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001100100000000000") port map( O =>C_59_S_2_L_4_out, I0 =>  inp_feat(493), I1 =>  inp_feat(440), I2 =>  inp_feat(112), I3 =>  inp_feat(22), I4 =>  inp_feat(51), I5 =>  inp_feat(11), I6 =>  inp_feat(341), I7 =>  inp_feat(219)); 
C_59_S_2_L_5_inst : LUT8 generic map(INIT => "0101010100000101000001010000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101100000001010100000000010100100000100000000001000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_2_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(362), I2 =>  inp_feat(158), I3 =>  inp_feat(358), I4 =>  inp_feat(45), I5 =>  inp_feat(400), I6 =>  inp_feat(89), I7 =>  inp_feat(177)); 
C_59_S_2_L_6_inst : LUT8 generic map(INIT => "1000101011000000000000000011111000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110010001100001011101000000000000000000000000000000000") port map( O =>C_59_S_2_L_6_out, I0 =>  inp_feat(431), I1 =>  inp_feat(66), I2 =>  inp_feat(473), I3 =>  inp_feat(476), I4 =>  inp_feat(412), I5 =>  inp_feat(277), I6 =>  inp_feat(507), I7 =>  inp_feat(397)); 
C_59_S_2_L_7_inst : LUT8 generic map(INIT => "0000010001110110000001110100011000000000000000000000000000000000000000100001101010000110000000100000000000001000000000000000001000010000011101001011011001000100000000000000000000000000000000000001000000110010010100100010000000000000000000000000000000000000") port map( O =>C_59_S_2_L_7_out, I0 =>  inp_feat(177), I1 =>  inp_feat(309), I2 =>  inp_feat(6), I3 =>  inp_feat(114), I4 =>  inp_feat(152), I5 =>  inp_feat(137), I6 =>  inp_feat(473), I7 =>  inp_feat(228)); 
C_59_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000100000000000000010000010000000001010101000001000000000101000000000000000000000000000001000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_3_L_0_out, I0 =>  inp_feat(359), I1 =>  inp_feat(271), I2 =>  inp_feat(238), I3 =>  inp_feat(288), I4 =>  inp_feat(418), I5 =>  inp_feat(4), I6 =>  inp_feat(441), I7 =>  inp_feat(277)); 
C_59_S_3_L_1_inst : LUT8 generic map(INIT => "0100011100000001000000010000000000011101010011010000000001001111000000000000000000000000000000000000000000000000000000000000000011101111000000101000000000000000111011110000101000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_3_L_1_out, I0 =>  inp_feat(218), I1 =>  inp_feat(221), I2 =>  inp_feat(416), I3 =>  inp_feat(91), I4 =>  inp_feat(408), I5 =>  inp_feat(182), I6 =>  inp_feat(277), I7 =>  inp_feat(441)); 
C_59_S_3_L_2_inst : LUT8 generic map(INIT => "0000000101000001000110001110000000000000000000000000000000000000010000000100000011111010111010000000000001001110001000000010011000000000001000000000000000110000000000000000000000000000000000000100000101000101100101100001100100000000000000000000000000000000") port map( O =>C_59_S_3_L_2_out, I0 =>  inp_feat(105), I1 =>  inp_feat(378), I2 =>  inp_feat(473), I3 =>  inp_feat(158), I4 =>  inp_feat(228), I5 =>  inp_feat(358), I6 =>  inp_feat(475), I7 =>  inp_feat(447)); 
C_59_S_3_L_3_inst : LUT8 generic map(INIT => "0000110000000000111010000000000010011101000010000000000000000000000001000000000000000000000000000101110101000100000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000100000000000000000000000000000") port map( O =>C_59_S_3_L_3_out, I0 =>  inp_feat(309), I1 =>  inp_feat(181), I2 =>  inp_feat(152), I3 =>  inp_feat(61), I4 =>  inp_feat(449), I5 =>  inp_feat(132), I6 =>  inp_feat(73), I7 =>  inp_feat(431)); 
C_59_S_3_L_4_inst : LUT8 generic map(INIT => "0000000001001100000000001110100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010001010111011001010111011111100100000000000000010000100000000010000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_3_L_4_out, I0 =>  inp_feat(45), I1 =>  inp_feat(400), I2 =>  inp_feat(47), I3 =>  inp_feat(158), I4 =>  inp_feat(362), I5 =>  inp_feat(270), I6 =>  inp_feat(89), I7 =>  inp_feat(177)); 
C_59_S_3_L_5_inst : LUT8 generic map(INIT => "0000001000000000101000100000000001010000000000000000101100000000001000001010000000100010000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_3_L_5_out, I0 =>  inp_feat(207), I1 =>  inp_feat(177), I2 =>  inp_feat(56), I3 =>  inp_feat(107), I4 =>  inp_feat(418), I5 =>  inp_feat(261), I6 =>  inp_feat(414), I7 =>  inp_feat(277)); 
C_59_S_3_L_6_inst : LUT8 generic map(INIT => "0000001000001001000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001010110000000000000011000000000000000000000000000000000000000000101000000000000000000000000000000000100000000000000011000000") port map( O =>C_59_S_3_L_6_out, I0 =>  inp_feat(223), I1 =>  inp_feat(210), I2 =>  inp_feat(437), I3 =>  inp_feat(497), I4 =>  inp_feat(66), I5 =>  inp_feat(358), I6 =>  inp_feat(385), I7 =>  inp_feat(261)); 
C_59_S_3_L_7_inst : LUT8 generic map(INIT => "0101000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000001010000000000000100000100000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_3_L_7_out, I0 =>  inp_feat(338), I1 =>  inp_feat(317), I2 =>  inp_feat(85), I3 =>  inp_feat(14), I4 =>  inp_feat(11), I5 =>  inp_feat(112), I6 =>  inp_feat(457), I7 =>  inp_feat(51)); 
C_59_S_4_L_0_inst : LUT8 generic map(INIT => "0000100000001000000010000000000000001000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000110000001000110000000000000000001100000000000000000000000000000010000000000000000000000000000000100000000000000000000000") port map( O =>C_59_S_4_L_0_out, I0 =>  inp_feat(494), I1 =>  inp_feat(14), I2 =>  inp_feat(317), I3 =>  inp_feat(507), I4 =>  inp_feat(245), I5 =>  inp_feat(426), I6 =>  inp_feat(69), I7 =>  inp_feat(182)); 
C_59_S_4_L_1_inst : LUT8 generic map(INIT => "1000000100010001001100001000011011000000100000000000000000000000000000000000000000000010000000001111001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000") port map( O =>C_59_S_4_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(399), I2 =>  inp_feat(274), I3 =>  inp_feat(396), I4 =>  inp_feat(352), I5 =>  inp_feat(476), I6 =>  inp_feat(228), I7 =>  inp_feat(431)); 
C_59_S_4_L_2_inst : LUT8 generic map(INIT => "0100100000000000000000000000000010001000000010000000000000000000000010001010110100000000100001000000000010001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000100010000000000000000000") port map( O =>C_59_S_4_L_2_out, I0 =>  inp_feat(101), I1 =>  inp_feat(50), I2 =>  inp_feat(184), I3 =>  inp_feat(41), I4 =>  inp_feat(224), I5 =>  inp_feat(75), I6 =>  inp_feat(341), I7 =>  inp_feat(219)); 
C_59_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010001000000000000000000000000000001000100000000000000000000000000010100000100010000010001010000011110001100100000000000000000000010100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000") port map( O =>C_59_S_4_L_3_out, I0 =>  inp_feat(488), I1 =>  inp_feat(51), I2 =>  inp_feat(411), I3 =>  inp_feat(101), I4 =>  inp_feat(471), I5 =>  inp_feat(184), I6 =>  inp_feat(198), I7 =>  inp_feat(4)); 
C_59_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000100011100100011100000000000000000000000000000010100000000000001111000100110011110100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000") port map( O =>C_59_S_4_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(87), I2 =>  inp_feat(322), I3 =>  inp_feat(130), I4 =>  inp_feat(418), I5 =>  inp_feat(329), I6 =>  inp_feat(483), I7 =>  inp_feat(457)); 
C_59_S_4_L_5_inst : LUT8 generic map(INIT => "0001000100101101001000000000101000000000000000000000000000000000000010001100111100101110000000000000000000000000001000000000000010100000000001011010000000000000000000000000000000100000000000001000000100000101000000000000000000000000000000001010000000000000") port map( O =>C_59_S_4_L_5_out, I0 =>  inp_feat(494), I1 =>  inp_feat(475), I2 =>  inp_feat(483), I3 =>  inp_feat(418), I4 =>  inp_feat(309), I5 =>  inp_feat(397), I6 =>  inp_feat(6), I7 =>  inp_feat(470)); 
C_59_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000001000000000000001000000000000110001000000000000000000000010001111110000000000110010100000000000101000000000000010000000000000100111010000000000000000000000000000000000000000000000000000000011010011000000000001111100000000000000000000000000000000") port map( O =>C_59_S_4_L_6_out, I0 =>  inp_feat(182), I1 =>  inp_feat(47), I2 =>  inp_feat(378), I3 =>  inp_feat(4), I4 =>  inp_feat(431), I5 =>  inp_feat(358), I6 =>  inp_feat(228), I7 =>  inp_feat(144)); 
C_59_S_4_L_7_inst : LUT8 generic map(INIT => "0111001000100000000001001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101000001000000000000000000110101111000010000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_59_S_4_L_7_out, I0 =>  inp_feat(41), I1 =>  inp_feat(75), I2 =>  inp_feat(391), I3 =>  inp_feat(507), I4 =>  inp_feat(223), I5 =>  inp_feat(55), I6 =>  inp_feat(457), I7 =>  inp_feat(470)); 
C_60_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110000000100001010001100100011000000010000000000000000000000000001000000000000000110000011000100000000000000000000000000100000") port map( O =>C_60_S_0_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(329), I2 =>  inp_feat(23), I3 =>  inp_feat(317), I4 =>  inp_feat(483), I5 =>  inp_feat(100), I6 =>  inp_feat(478), I7 =>  inp_feat(488)); 
C_60_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001100000000000000000000000000000000000000000000001100000000000000111000001010000000000000000000000000000010000000") port map( O =>C_60_S_0_L_1_out, I0 =>  inp_feat(504), I1 =>  inp_feat(285), I2 =>  inp_feat(408), I3 =>  inp_feat(396), I4 =>  inp_feat(483), I5 =>  inp_feat(445), I6 =>  inp_feat(108), I7 =>  inp_feat(226)); 
C_60_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000001000000000000000000000001000000100000000000000000000000000001000000000000000000010000000100010001000000010000000000000000000000110000000000000001001000010000001000000011000000000000000100010111010000010000000000000001000000010000000100") port map( O =>C_60_S_0_L_2_out, I0 =>  inp_feat(483), I1 =>  inp_feat(143), I2 =>  inp_feat(488), I3 =>  inp_feat(494), I4 =>  inp_feat(318), I5 =>  inp_feat(335), I6 =>  inp_feat(152), I7 =>  inp_feat(407)); 
C_60_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000000000001000000000101100010011001000000000000100000010000100010001001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_0_L_3_out, I0 =>  inp_feat(317), I1 =>  inp_feat(329), I2 =>  inp_feat(387), I3 =>  inp_feat(196), I4 =>  inp_feat(269), I5 =>  inp_feat(251), I6 =>  inp_feat(483), I7 =>  inp_feat(408)); 
C_60_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000010001010000000000000100010001000101010101010101010000000000000000000000000000010001100000000001100000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000") port map( O =>C_60_S_0_L_4_out, I0 =>  inp_feat(436), I1 =>  inp_feat(441), I2 =>  inp_feat(182), I3 =>  inp_feat(114), I4 =>  inp_feat(308), I5 =>  inp_feat(483), I6 =>  inp_feat(265), I7 =>  inp_feat(100)); 
C_60_S_0_L_5_inst : LUT8 generic map(INIT => "0011000100000000000000000000000001110101000011000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010100000100010000000000000000000000000000000100000001000000000000000100010001000100000000000000") port map( O =>C_60_S_0_L_5_out, I0 =>  inp_feat(488), I1 =>  inp_feat(476), I2 =>  inp_feat(294), I3 =>  inp_feat(73), I4 =>  inp_feat(130), I5 =>  inp_feat(483), I6 =>  inp_feat(94), I7 =>  inp_feat(256)); 
C_60_S_0_L_6_inst : LUT8 generic map(INIT => "0000010000000100000001001100010000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000001010001000101010001000100000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_0_L_6_out, I0 =>  inp_feat(488), I1 =>  inp_feat(190), I2 =>  inp_feat(172), I3 =>  inp_feat(114), I4 =>  inp_feat(152), I5 =>  inp_feat(304), I6 =>  inp_feat(408), I7 =>  inp_feat(218)); 
C_60_S_0_L_7_inst : LUT8 generic map(INIT => "0000011100000000000101010000000000000000000000000000000000000100011001010000000011000101000000000000000000000000000000000000000000000000000001010000010000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000") port map( O =>C_60_S_0_L_7_out, I0 =>  inp_feat(488), I1 =>  inp_feat(504), I2 =>  inp_feat(187), I3 =>  inp_feat(254), I4 =>  inp_feat(475), I5 =>  inp_feat(143), I6 =>  inp_feat(238), I7 =>  inp_feat(256)); 
C_60_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110000000100001010001100100011000000010000000000000000000000000001000000000000000110000011000100000000000000000000000000100000") port map( O =>C_60_S_1_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(329), I2 =>  inp_feat(23), I3 =>  inp_feat(317), I4 =>  inp_feat(483), I5 =>  inp_feat(100), I6 =>  inp_feat(478), I7 =>  inp_feat(488)); 
C_60_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001000100100000000000000000000000000000000000000010000100000000000000000000010001000000000000000000000000000000000000000000000000000100010000000001000100000000000000010000000000000001000000000000010111100001011") port map( O =>C_60_S_1_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(152), I2 =>  inp_feat(488), I3 =>  inp_feat(376), I4 =>  inp_feat(283), I5 =>  inp_feat(483), I6 =>  inp_feat(108), I7 =>  inp_feat(226)); 
C_60_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000010000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001010100000101000000000000010000000000010001000000000000000000000000000000010000000000000000000000000000000000000000000001010100000101000001010") port map( O =>C_60_S_1_L_2_out, I0 =>  inp_feat(408), I1 =>  inp_feat(347), I2 =>  inp_feat(483), I3 =>  inp_feat(318), I4 =>  inp_feat(308), I5 =>  inp_feat(204), I6 =>  inp_feat(476), I7 =>  inp_feat(187)); 
C_60_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000100000000000000000000000000000000000000000011001111100011001000110000001100000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000000000000010000000000000000000000") port map( O =>C_60_S_1_L_3_out, I0 =>  inp_feat(251), I1 =>  inp_feat(190), I2 =>  inp_feat(207), I3 =>  inp_feat(222), I4 =>  inp_feat(441), I5 =>  inp_feat(32), I6 =>  inp_feat(488), I7 =>  inp_feat(304)); 
C_60_S_1_L_4_inst : LUT8 generic map(INIT => "0100000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000011111110001010100000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000") port map( O =>C_60_S_1_L_4_out, I0 =>  inp_feat(437), I1 =>  inp_feat(399), I2 =>  inp_feat(265), I3 =>  inp_feat(60), I4 =>  inp_feat(61), I5 =>  inp_feat(493), I6 =>  inp_feat(190), I7 =>  inp_feat(483)); 
C_60_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000001000000010100000111000001100000011000000000000000000000000000000000000000000000000110000000000000000000000000000001000000000000000000000000000001100000000000000000000000000000000100000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_1_L_5_out, I0 =>  inp_feat(304), I1 =>  inp_feat(269), I2 =>  inp_feat(408), I3 =>  inp_feat(251), I4 =>  inp_feat(335), I5 =>  inp_feat(483), I6 =>  inp_feat(190), I7 =>  inp_feat(242)); 
C_60_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000010000000000000011000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000011000000100010000000000000000000110000001100100011000000010000000000000000000000000000000000000001000000100010000000000000000000") port map( O =>C_60_S_1_L_6_out, I0 =>  inp_feat(494), I1 =>  inp_feat(493), I2 =>  inp_feat(436), I3 =>  inp_feat(170), I4 =>  inp_feat(78), I5 =>  inp_feat(152), I6 =>  inp_feat(478), I7 =>  inp_feat(318)); 
C_60_S_1_L_7_inst : LUT8 generic map(INIT => "1000000000001101000010000001010000000000000001000001000001010000000000000000000000000000010000000000000000000000000000000000000000001100100011000000000000000100000000000000010000010001000001010000000000000000000000000000000000000000000000000101000001000000") port map( O =>C_60_S_1_L_7_out, I0 =>  inp_feat(310), I1 =>  inp_feat(478), I2 =>  inp_feat(226), I3 =>  inp_feat(152), I4 =>  inp_feat(98), I5 =>  inp_feat(256), I6 =>  inp_feat(242), I7 =>  inp_feat(29)); 
C_60_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110000000100001010001100100011000000010000000000000000000000000001000000000000000110000011000100000000000000000000000000100000") port map( O =>C_60_S_2_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(329), I2 =>  inp_feat(23), I3 =>  inp_feat(317), I4 =>  inp_feat(483), I5 =>  inp_feat(100), I6 =>  inp_feat(478), I7 =>  inp_feat(488)); 
C_60_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001000100100000000000000000000000000000000000000010000100000000000000000000010001000000000000000000000000000000000000000000000000000100010000000001000100000000000000010000000000000001000000000000010111100001011") port map( O =>C_60_S_2_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(152), I2 =>  inp_feat(488), I3 =>  inp_feat(376), I4 =>  inp_feat(283), I5 =>  inp_feat(483), I6 =>  inp_feat(108), I7 =>  inp_feat(226)); 
C_60_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000010000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001010100000101000000000000010000000000010001000000000000000000000000000000010000000000000000000000000000000000000000000001010100000101000001010") port map( O =>C_60_S_2_L_2_out, I0 =>  inp_feat(408), I1 =>  inp_feat(347), I2 =>  inp_feat(483), I3 =>  inp_feat(318), I4 =>  inp_feat(308), I5 =>  inp_feat(204), I6 =>  inp_feat(476), I7 =>  inp_feat(187)); 
C_60_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000100000000000000000000000000000000000000000011001111100011001000110000001100000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000000000000010000000000000000000000") port map( O =>C_60_S_2_L_3_out, I0 =>  inp_feat(251), I1 =>  inp_feat(190), I2 =>  inp_feat(207), I3 =>  inp_feat(222), I4 =>  inp_feat(441), I5 =>  inp_feat(32), I6 =>  inp_feat(488), I7 =>  inp_feat(304)); 
C_60_S_2_L_4_inst : LUT8 generic map(INIT => "0000100000001000000000001000100000000000101000000000000000000000100010001010100010101000101010001000100010100000101010000010000000000000000000000000000000000000000000000100000000000000000000000001100000010000000000000111000000000000101000000010000010000000") port map( O =>C_60_S_2_L_4_out, I0 =>  inp_feat(190), I1 =>  inp_feat(317), I2 =>  inp_feat(115), I3 =>  inp_feat(182), I4 =>  inp_feat(221), I5 =>  inp_feat(256), I6 =>  inp_feat(483), I7 =>  inp_feat(478)); 
C_60_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000001000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010001100011001100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_2_L_5_out, I0 =>  inp_feat(416), I1 =>  inp_feat(157), I2 =>  inp_feat(434), I3 =>  inp_feat(251), I4 =>  inp_feat(335), I5 =>  inp_feat(61), I6 =>  inp_feat(493), I7 =>  inp_feat(483)); 
C_60_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000010000000000000001100000100000000000000000000000000000000100000000010000010100001101000001010000010100000101000000100000000000000010000000000000101000001000000000100000001000000000000000000000000000000000000001000000010000000001000000000000") port map( O =>C_60_S_2_L_6_out, I0 =>  inp_feat(476), I1 =>  inp_feat(83), I2 =>  inp_feat(61), I3 =>  inp_feat(221), I4 =>  inp_feat(201), I5 =>  inp_feat(483), I6 =>  inp_feat(418), I7 =>  inp_feat(256)); 
C_60_S_2_L_7_inst : LUT8 generic map(INIT => "0000000100000000000001000000000000000110000010000000110100000000000000000000000001000100000000000000010000000000000011010000000001000000000000000000100000000000000011010000000000001111000000001000000000001010100011000000100000001111000001000000110110000001") port map( O =>C_60_S_2_L_7_out, I0 =>  inp_feat(375), I1 =>  inp_feat(16), I2 =>  inp_feat(483), I3 =>  inp_feat(130), I4 =>  inp_feat(416), I5 =>  inp_feat(152), I6 =>  inp_feat(29), I7 =>  inp_feat(308)); 
C_60_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110000000100001010001100100011000000010000000000000000000000000001000000000000000110000011000100000000000000000000000000100000") port map( O =>C_60_S_3_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(329), I2 =>  inp_feat(23), I3 =>  inp_feat(317), I4 =>  inp_feat(483), I5 =>  inp_feat(100), I6 =>  inp_feat(478), I7 =>  inp_feat(488)); 
C_60_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001000100100000000000000000000000000000000000000010000100000000000000000000010001000000000000000000000000000000000000000000000000000100010000000001000100000000000000010000000000000001000000000000010111100001011") port map( O =>C_60_S_3_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(152), I2 =>  inp_feat(488), I3 =>  inp_feat(376), I4 =>  inp_feat(283), I5 =>  inp_feat(483), I6 =>  inp_feat(108), I7 =>  inp_feat(226)); 
C_60_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100000110000000000000000001000000000000100000000000000000000000000000000000000100000000000000000000010010000010000000011000110110001001100000000000000000000000000001011000000000000000000000000") port map( O =>C_60_S_3_L_2_out, I0 =>  inp_feat(152), I1 =>  inp_feat(483), I2 =>  inp_feat(488), I3 =>  inp_feat(265), I4 =>  inp_feat(317), I5 =>  inp_feat(336), I6 =>  inp_feat(476), I7 =>  inp_feat(187)); 
C_60_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000010000000000000000000000010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000001000000000101000100010001000000000000010110000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_3_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(483), I2 =>  inp_feat(318), I3 =>  inp_feat(336), I4 =>  inp_feat(434), I5 =>  inp_feat(251), I6 =>  inp_feat(493), I7 =>  inp_feat(467)); 
C_60_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000100000001001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010110000011100001100000011010000101000000001000000000000101100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_3_L_4_out, I0 =>  inp_feat(73), I1 =>  inp_feat(256), I2 =>  inp_feat(136), I3 =>  inp_feat(328), I4 =>  inp_feat(251), I5 =>  inp_feat(23), I6 =>  inp_feat(332), I7 =>  inp_feat(483)); 
C_60_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000011000010000000000000000000000000001000100000000000000000010000000000000000000000000000000000000000000010000000000000000010000000010000100000000000000010000000000010001010000000000000111100001000000000000000000000000000000000000000100000000000") port map( O =>C_60_S_3_L_5_out, I0 =>  inp_feat(94), I1 =>  inp_feat(256), I2 =>  inp_feat(488), I3 =>  inp_feat(352), I4 =>  inp_feat(437), I5 =>  inp_feat(441), I6 =>  inp_feat(294), I7 =>  inp_feat(475)); 
C_60_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000101000100001100100100000000000000000000001000101010000000000000000001000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000100000001000000000000000000000000000000000") port map( O =>C_60_S_3_L_6_out, I0 =>  inp_feat(204), I1 =>  inp_feat(91), I2 =>  inp_feat(182), I3 =>  inp_feat(488), I4 =>  inp_feat(483), I5 =>  inp_feat(317), I6 =>  inp_feat(378), I7 =>  inp_feat(445)); 
C_60_S_3_L_7_inst : LUT8 generic map(INIT => "0100010001001100000001000000110111010100000001000000000000000000000000000000000000000000000000000000010000000000000001010000000100000000000000000000010000000101000001000000000000000000000011000000000000000000000000000000000000000000000000000000000000000101") port map( O =>C_60_S_3_L_7_out, I0 =>  inp_feat(483), I1 =>  inp_feat(478), I2 =>  inp_feat(318), I3 =>  inp_feat(182), I4 =>  inp_feat(379), I5 =>  inp_feat(475), I6 =>  inp_feat(195), I7 =>  inp_feat(23)); 
C_60_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110000000100001010001100100011000000010000000000000000000000000001000000000000000110000011000100000000000000000000000000100000") port map( O =>C_60_S_4_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(329), I2 =>  inp_feat(23), I3 =>  inp_feat(317), I4 =>  inp_feat(483), I5 =>  inp_feat(100), I6 =>  inp_feat(478), I7 =>  inp_feat(488)); 
C_60_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000001000100100000000000000000000000000000000000000010000100000000000000000000010001000000000000000000000000000000000000000000000000000100010000000001000100000000000000010000000000000001000000000000010111100001011") port map( O =>C_60_S_4_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(152), I2 =>  inp_feat(488), I3 =>  inp_feat(376), I4 =>  inp_feat(283), I5 =>  inp_feat(483), I6 =>  inp_feat(108), I7 =>  inp_feat(226)); 
C_60_S_4_L_2_inst : LUT8 generic map(INIT => "0000000001000000000000000100000000000000010001000000000001000000000000000000010010000000010000000100000001000000000000001100000000000000000000000000000000000000010000001111010100000000010000000000000000000000000000000100000000000000100000000000000011000000") port map( O =>C_60_S_4_L_2_out, I0 =>  inp_feat(483), I1 =>  inp_feat(190), I2 =>  inp_feat(23), I3 =>  inp_feat(488), I4 =>  inp_feat(494), I5 =>  inp_feat(318), I6 =>  inp_feat(441), I7 =>  inp_feat(294)); 
C_60_S_4_L_3_inst : LUT8 generic map(INIT => "0010111000101010000000000010101000000000000010000011111100100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_4_L_3_out, I0 =>  inp_feat(478), I1 =>  inp_feat(251), I2 =>  inp_feat(483), I3 =>  inp_feat(114), I4 =>  inp_feat(294), I5 =>  inp_feat(212), I6 =>  inp_feat(136), I7 =>  inp_feat(408)); 
C_60_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000010000000000000000000000000000000000000100011111010100000000000100000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000001000000010100000000000001000000000000000000000000000000000000000") port map( O =>C_60_S_4_L_4_out, I0 =>  inp_feat(297), I1 =>  inp_feat(256), I2 =>  inp_feat(269), I3 =>  inp_feat(483), I4 =>  inp_feat(304), I5 =>  inp_feat(408), I6 =>  inp_feat(488), I7 =>  inp_feat(476)); 
C_60_S_4_L_5_inst : LUT8 generic map(INIT => "0010000000000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_60_S_4_L_5_out, I0 =>  inp_feat(100), I1 =>  inp_feat(182), I2 =>  inp_feat(493), I3 =>  inp_feat(332), I4 =>  inp_feat(61), I5 =>  inp_feat(152), I6 =>  inp_feat(305), I7 =>  inp_feat(476)); 
C_60_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000001010000000000000000000000000000010000000000000000000000010001101110000000000000000000000000011001100000000000000000000000000000010000000000000000000000010000000100000000000000000000000000000101000000000000000000001000000011110000000000000000000") port map( O =>C_60_S_4_L_6_out, I0 =>  inp_feat(256), I1 =>  inp_feat(317), I2 =>  inp_feat(476), I3 =>  inp_feat(483), I4 =>  inp_feat(61), I5 =>  inp_feat(182), I6 =>  inp_feat(301), I7 =>  inp_feat(328)); 
C_60_S_4_L_7_inst : LUT8 generic map(INIT => "0000010100001101010110011101010100000000000000000001000000000000000000000000000000010011000000000000000000000000010100000000000000000000000000010000010100000000000000000000000000010000000000000000000000000100000001010000000000000000000000000000000000000000") port map( O =>C_60_S_4_L_7_out, I0 =>  inp_feat(483), I1 =>  inp_feat(152), I2 =>  inp_feat(308), I3 =>  inp_feat(441), I4 =>  inp_feat(318), I5 =>  inp_feat(436), I6 =>  inp_feat(23), I7 =>  inp_feat(478)); 
C_61_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_0_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_1_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_2_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_3_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_0_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_1_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_2_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_3_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_4_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_5_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_6_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_61_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000") port map( O =>C_61_S_4_L_7_out, I0 =>  inp_feat(3), I1 =>  inp_feat(2), I2 =>  inp_feat(1), I3 =>  inp_feat(0), I4 =>  inp_feat(50), I5 =>  inp_feat(204), I6 =>  inp_feat(418), I7 =>  inp_feat(488)); 
C_62_S_0_L_0_inst : LUT8 generic map(INIT => "1111110111111111110011001111110111111101111101011111010011110101101000001100110110100000000001011111000001110101101000001111010100000000101000000000000000010000010100000001000100000000111100000000000000001000000000000000000000000000000000000000000000010001") port map( O =>C_62_S_0_L_0_out, I0 =>  inp_feat(100), I1 =>  inp_feat(6), I2 =>  inp_feat(416), I3 =>  inp_feat(98), I4 =>  inp_feat(431), I5 =>  inp_feat(190), I6 =>  inp_feat(187), I7 =>  inp_feat(488)); 
C_62_S_0_L_1_inst : LUT8 generic map(INIT => "1110000011001000110000001000000011111010000000001110000010000000010000000000000000000000100000001111000010100000101000001000000011100100110000001100000001000000111111111110111011100000100000000100000000000000000000000000000011000011010001001010000010001000") port map( O =>C_62_S_0_L_1_out, I0 =>  inp_feat(493), I1 =>  inp_feat(139), I2 =>  inp_feat(488), I3 =>  inp_feat(483), I4 =>  inp_feat(449), I5 =>  inp_feat(461), I6 =>  inp_feat(380), I7 =>  inp_feat(365)); 
C_62_S_0_L_2_inst : LUT8 generic map(INIT => "1111111111110101101000001011000100110000110101001000000010010000001000011011000010100000001000000000000000100000101000010111000011111101011101011000000100010001110111000101000010000001010100001010110000100000101011111111011110000000000000001000101101010000") port map( O =>C_62_S_0_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(61), I2 =>  inp_feat(256), I3 =>  inp_feat(107), I4 =>  inp_feat(232), I5 =>  inp_feat(504), I6 =>  inp_feat(407), I7 =>  inp_feat(457)); 
C_62_S_0_L_3_inst : LUT8 generic map(INIT => "1111110011101000110100001000000011110000101000000001000010000000001000001010100000000000000000001100000010100000000000000000000011111000000000000100000000000000010100000000000000000000000000001101000000000000000000000000000011110000000000000000000000000000") port map( O =>C_62_S_0_L_3_out, I0 =>  inp_feat(221), I1 =>  inp_feat(91), I2 =>  inp_feat(446), I3 =>  inp_feat(359), I4 =>  inp_feat(418), I5 =>  inp_feat(504), I6 =>  inp_feat(407), I7 =>  inp_feat(37)); 
C_62_S_0_L_4_inst : LUT8 generic map(INIT => "1111101011111110101000101010001010101010110011000000001011101100111111101000000011000000100000000010001000000000000000000000000010101011000100001010000000000000011011100000000000000000000000000010001000000000000000000000000000000000000000000000000000000000") port map( O =>C_62_S_0_L_4_out, I0 =>  inp_feat(187), I1 =>  inp_feat(100), I2 =>  inp_feat(355), I3 =>  inp_feat(288), I4 =>  inp_feat(418), I5 =>  inp_feat(476), I6 =>  inp_feat(275), I7 =>  inp_feat(182)); 
C_62_S_0_L_5_inst : LUT8 generic map(INIT => "1110110000101010110011101010111011000000000010101100000001001010100100000000000011101100000011000000000000000000110010000101110011101000101001001010110011101111000000000000000000000100010010110000000000000000101011001100110000000000000001000000000001001101") port map( O =>C_62_S_0_L_5_out, I0 =>  inp_feat(139), I1 =>  inp_feat(483), I2 =>  inp_feat(318), I3 =>  inp_feat(407), I4 =>  inp_feat(478), I5 =>  inp_feat(182), I6 =>  inp_feat(403), I7 =>  inp_feat(457)); 
C_62_S_0_L_6_inst : LUT8 generic map(INIT => "0111111101101110001111010000001011001101110011010100110001000000111100010011011100000100010001010100010101010101010001000000010011111111111101111010000010000000110101011101010101000100000000011110000111111111000000000001000001000101111111010100000000000000") port map( O =>C_62_S_0_L_6_out, I0 =>  inp_feat(61), I1 =>  inp_feat(23), I2 =>  inp_feat(493), I3 =>  inp_feat(306), I4 =>  inp_feat(152), I5 =>  inp_feat(244), I6 =>  inp_feat(403), I7 =>  inp_feat(457)); 
C_62_S_0_L_7_inst : LUT8 generic map(INIT => "1101111111111101010100111101111111111111110100010011001101010001101100100111000100000101111000010111111111110111001100111111001101001001011101110001001101010001111100111101000100110011010100010000010000010000000000010000000000100011011100000011001101010001") port map( O =>C_62_S_0_L_7_out, I0 =>  inp_feat(408), I1 =>  inp_feat(143), I2 =>  inp_feat(304), I3 =>  inp_feat(201), I4 =>  inp_feat(174), I5 =>  inp_feat(195), I6 =>  inp_feat(222), I7 =>  inp_feat(472)); 
C_62_S_1_L_0_inst : LUT8 generic map(INIT => "1111110011011000111111101100000011100000000000000010000000000000111101010100000000000000000000001010000000000000000000000000000111110111010100000111100011000000111111111111011111100111111100101111010111001100111110001110010011101111111111111111111111111111") port map( O =>C_62_S_1_L_0_out, I0 =>  inp_feat(265), I1 =>  inp_feat(87), I2 =>  inp_feat(79), I3 =>  inp_feat(137), I4 =>  inp_feat(472), I5 =>  inp_feat(242), I6 =>  inp_feat(403), I7 =>  inp_feat(365)); 
C_62_S_1_L_1_inst : LUT8 generic map(INIT => "1110111111111111111011101110110000001100110011001010101011101000101011110000101100100000000000000000000001000000001000000000000011001100010111000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000") port map( O =>C_62_S_1_L_1_out, I0 =>  inp_feat(222), I1 =>  inp_feat(69), I2 =>  inp_feat(107), I3 =>  inp_feat(323), I4 =>  inp_feat(209), I5 =>  inp_feat(437), I6 =>  inp_feat(283), I7 =>  inp_feat(488)); 
C_62_S_1_L_2_inst : LUT8 generic map(INIT => "1011111011101111110010001000000101101000101010001010001010001010011000011100001100000001111000110000000000001010000000000000000011101110000011111100111110001011100010000000001000000000000010101011101100001011101010111010101100000000000010000000000000001010") port map( O =>C_62_S_1_L_2_out, I0 =>  inp_feat(475), I1 =>  inp_feat(493), I2 =>  inp_feat(218), I3 =>  inp_feat(207), I4 =>  inp_feat(387), I5 =>  inp_feat(483), I6 =>  inp_feat(283), I7 =>  inp_feat(61)); 
C_62_S_1_L_3_inst : LUT8 generic map(INIT => "1111111110101000111010001010101000000000000000000000000000000000111100101011001010100000101000100000000000000000000000000000000010111010101010101011111110011010000000011110000000010000000000001101000100011000001100000011000000010000001000000000000100100000") port map( O =>C_62_S_1_L_3_out, I0 =>  inp_feat(483), I1 =>  inp_feat(408), I2 =>  inp_feat(91), I3 =>  inp_feat(265), I4 =>  inp_feat(69), I5 =>  inp_feat(488), I6 =>  inp_feat(87), I7 =>  inp_feat(218)); 
C_62_S_1_L_4_inst : LUT8 generic map(INIT => "0110101110100000111110000000100011111000000000001010100000000000000000000000100011001010000010001000000000000000101000000000000001101111101110001111111111111110010100000000000001000000000000000000011000001000101010011110111100000000000000000000000000000000") port map( O =>C_62_S_1_L_4_out, I0 =>  inp_feat(87), I1 =>  inp_feat(460), I2 =>  inp_feat(195), I3 =>  inp_feat(304), I4 =>  inp_feat(100), I5 =>  inp_feat(345), I6 =>  inp_feat(182), I7 =>  inp_feat(478)); 
C_62_S_1_L_5_inst : LUT8 generic map(INIT => "1110100011100000110010001111000011110000100000000000000010000000100010001000000011001000100000001110000010000000110000001000000011101010110010101100110010110000100000001100110011001000110110001000000000000000110000000000000010000000000000001000000000000000") port map( O =>C_62_S_1_L_5_out, I0 =>  inp_feat(483), I1 =>  inp_feat(459), I2 =>  inp_feat(329), I3 =>  inp_feat(336), I4 =>  inp_feat(379), I5 =>  inp_feat(79), I6 =>  inp_feat(345), I7 =>  inp_feat(478)); 
C_62_S_1_L_6_inst : LUT8 generic map(INIT => "1110111000000000001010000000100011001100000000000000100000001000101010001000100010101000000010001000100000000000100010001010100011101010110010000000000000000000000000000000000000001000000000001100101100001110101000000000000010001000000000000000100000000000") port map( O =>C_62_S_1_L_6_out, I0 =>  inp_feat(210), I1 =>  inp_feat(271), I2 =>  inp_feat(288), I3 =>  inp_feat(476), I4 =>  inp_feat(40), I5 =>  inp_feat(329), I6 =>  inp_feat(478), I7 =>  inp_feat(336)); 
C_62_S_1_L_7_inst : LUT8 generic map(INIT => "1110110011100000100000000000000011010101000000001110110100000000110000001110000000000100000000000000000000000000000000000000000011111100110101001100010001000000110001001100000011001000000000001000010011000000110001000000000010000000000000001000000000000000") port map( O =>C_62_S_1_L_7_out, I0 =>  inp_feat(474), I1 =>  inp_feat(418), I2 =>  inp_feat(459), I3 =>  inp_feat(329), I4 =>  inp_feat(483), I5 =>  inp_feat(51), I6 =>  inp_feat(91), I7 =>  inp_feat(190)); 
C_62_S_2_L_0_inst : LUT8 generic map(INIT => "1010111010001000100011110000000111101110100010000000111000000000100011001010101000001110000010101010111110101110001011100000101010001110100000001000101000101000100010000011100000000000000000100010101000101010001010100010101110101010001010000000101000100011") port map( O =>C_62_S_2_L_0_out, I0 =>  inp_feat(488), I1 =>  inp_feat(128), I2 =>  inp_feat(190), I3 =>  inp_feat(342), I4 =>  inp_feat(182), I5 =>  inp_feat(229), I6 =>  inp_feat(457), I7 =>  inp_feat(187)); 
C_62_S_2_L_1_inst : LUT8 generic map(INIT => "1111110011000000111111001100010000001000000010001111100011010100111110001100000011000001010101011000100000000000001100011111110111110000110011000111010011001101000001000000000001000000100000011000100111001101100101011101010110001111100011111111010000110111") port map( O =>C_62_S_2_L_1_out, I0 =>  inp_feat(408), I1 =>  inp_feat(403), I2 =>  inp_feat(269), I3 =>  inp_feat(60), I4 =>  inp_feat(436), I5 =>  inp_feat(187), I6 =>  inp_feat(61), I7 =>  inp_feat(218)); 
C_62_S_2_L_2_inst : LUT8 generic map(INIT => "1101111011010100111011111100111111111100110111000100010001000100111010001100000010001110000000000100000000000000000001000000000011010000110100011100110111001111110010001101010011000001110011001101010111010000000001000100010111000100010101000000010001000101") port map( O =>C_62_S_2_L_2_out, I0 =>  inp_feat(100), I1 =>  inp_feat(483), I2 =>  inp_feat(306), I3 =>  inp_feat(411), I4 =>  inp_feat(387), I5 =>  inp_feat(132), I6 =>  inp_feat(69), I7 =>  inp_feat(81)); 
C_62_S_2_L_3_inst : LUT8 generic map(INIT => "1111111011001100100000101100100011101111110011110000100010101010010011000100110010000000000000000100100111011111000010000000000011111111110011111011100011001000000001111000111100000000001010001100110011001111000000001100001010001000001011100000000010001010") port map( O =>C_62_S_2_L_3_out, I0 =>  inp_feat(469), I1 =>  inp_feat(172), I2 =>  inp_feat(190), I3 =>  inp_feat(137), I4 =>  inp_feat(489), I5 =>  inp_feat(6), I6 =>  inp_feat(318), I7 =>  inp_feat(221)); 
C_62_S_2_L_4_inst : LUT8 generic map(INIT => "1010111011100110000011000001000011111101110111001101000111010101111011100010001011100111001100011111110111110101111101111111011111000000110011000000000000000000110000001100110101000100010100000000000000000000000001000000000000010001010101010000000001010101") port map( O =>C_62_S_2_L_4_out, I0 =>  inp_feat(81), I1 =>  inp_feat(290), I2 =>  inp_feat(265), I3 =>  inp_feat(497), I4 =>  inp_feat(251), I5 =>  inp_feat(61), I6 =>  inp_feat(242), I7 =>  inp_feat(91)); 
C_62_S_2_L_5_inst : LUT8 generic map(INIT => "1111001010001010000000110000101010000000100000000000000000000000111111110001101001011111011100101100000000000000000101000111001011111011001110110010001100101000100000000000000100000000000000001111111101111110011111110111111111011100010000000101010001010100") port map( O =>C_62_S_2_L_5_out, I0 =>  inp_feat(445), I1 =>  inp_feat(242), I2 =>  inp_feat(444), I3 =>  inp_feat(265), I4 =>  inp_feat(403), I5 =>  inp_feat(91), I6 =>  inp_feat(61), I7 =>  inp_feat(408)); 
C_62_S_2_L_6_inst : LUT8 generic map(INIT => "0100010011111101111110111101010111010001111111010111111011110110110100000100000011000000000000001001000010000000000100000000000001000100111011001101000101010001100101001100010000000001011101011100110011000000110011000000000011110000011100000111000001010000") port map( O =>C_62_S_2_L_6_out, I0 =>  inp_feat(408), I1 =>  inp_feat(60), I2 =>  inp_feat(218), I3 =>  inp_feat(291), I4 =>  inp_feat(143), I5 =>  inp_feat(398), I6 =>  inp_feat(175), I7 =>  inp_feat(114)); 
C_62_S_2_L_7_inst : LUT8 generic map(INIT => "1111000001111000011000001010000011010000111100001001100000000000011100000000000000010010000000000001000110101000101110110000100011100000000000001111100000000000101100000010000011111000001000001101000000000000001000000010000011100000110011101111100000011001") port map( O =>C_62_S_2_L_7_out, I0 =>  inp_feat(256), I1 =>  inp_feat(172), I2 =>  inp_feat(488), I3 =>  inp_feat(483), I4 =>  inp_feat(322), I5 =>  inp_feat(195), I6 =>  inp_feat(222), I7 =>  inp_feat(61)); 
C_62_S_3_L_0_inst : LUT8 generic map(INIT => "1111101011111111111000000010001011100011001000000001001000100000111000000010001000100000001000001001100111111100101000100010000010101010101011111000000010000000111000101111001000000000000000001010100010101010000000000000000011110011111100100000000000000000") port map( O =>C_62_S_3_L_0_out, I0 =>  inp_feat(304), I1 =>  inp_feat(408), I2 =>  inp_feat(483), I3 =>  inp_feat(290), I4 =>  inp_feat(459), I5 =>  inp_feat(468), I6 =>  inp_feat(37), I7 =>  inp_feat(457)); 
C_62_S_3_L_1_inst : LUT8 generic map(INIT => "0101101010101000111101011111110100101111100011001101110100000001101110111110100011011101111111011011111110001000010111110101010101010111011000010001010111010111010111000000000011000101000001111000000000000000000011010001110110001100000110100001110100011101") port map( O =>C_62_S_3_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(79), I2 =>  inp_feat(190), I3 =>  inp_feat(291), I4 =>  inp_feat(457), I5 =>  inp_feat(6), I6 =>  inp_feat(37), I7 =>  inp_feat(336)); 
C_62_S_3_L_2_inst : LUT8 generic map(INIT => "1111111111001110110100011000000010000000000010001100010100000000111011101000001011001001000000001110110010101000110011000000000011111111011011101000110010101010000000000000000000000000000000001001111110000011000000000000000000000000000000000000000000000000") port map( O =>C_62_S_3_L_2_out, I0 =>  inp_feat(416), I1 =>  inp_feat(317), I2 =>  inp_feat(408), I3 =>  inp_feat(222), I4 =>  inp_feat(359), I5 =>  inp_feat(504), I6 =>  inp_feat(472), I7 =>  inp_feat(444)); 
C_62_S_3_L_3_inst : LUT8 generic map(INIT => "0111101010111010111111111110010100111101000100000010001111011011100111101111001010101011011000100000001000000000000000011101100011011111100110101011101111111111000111110000100000111111011111111011111110110110101111111111111100001001000100000010111110110111") port map( O =>C_62_S_3_L_3_out, I0 =>  inp_feat(472), I1 =>  inp_feat(408), I2 =>  inp_feat(221), I3 =>  inp_feat(87), I4 =>  inp_feat(387), I5 =>  inp_feat(342), I6 =>  inp_feat(229), I7 =>  inp_feat(457)); 
C_62_S_3_L_4_inst : LUT8 generic map(INIT => "1101100011001000110111001100110011001100010000001000110001000100110010000100000011010100010001001101110001000000110101000100000010101010101000000000010011100100000000001100000000000100011000001000000001000000110001000100010000001000000000001100110001000100") port map( O =>C_62_S_3_L_4_out, I0 =>  inp_feat(413), I1 =>  inp_feat(476), I2 =>  inp_feat(380), I3 =>  inp_feat(51), I4 =>  inp_feat(100), I5 =>  inp_feat(130), I6 =>  inp_feat(465), I7 =>  inp_feat(328)); 
C_62_S_3_L_5_inst : LUT8 generic map(INIT => "1101011101101111011100111100010001011111001101010001010101000010011011000010000000100000001011000101010100000001000001110000010111011111010001011101000111000100010001010001111100010101010101011000010000000000000000000000000001000101000001000000000001000000") port map( O =>C_62_S_3_L_5_out, I0 =>  inp_feat(61), I1 =>  inp_feat(23), I2 =>  inp_feat(143), I3 =>  inp_feat(130), I4 =>  inp_feat(29), I5 =>  inp_feat(445), I6 =>  inp_feat(152), I7 =>  inp_feat(244)); 
C_62_S_3_L_6_inst : LUT8 generic map(INIT => "0010111000011110111111000110110011001100000010000100110001011101000010101010101001001000100011001000100010000000010010000100000101011110010111110000010000001100000010000000110000000000000001000010101000101110000000000000110000001000100011100000000001001110") port map( O =>C_62_S_3_L_6_out, I0 =>  inp_feat(221), I1 =>  inp_feat(152), I2 =>  inp_feat(100), I3 =>  inp_feat(73), I4 =>  inp_feat(387), I5 =>  inp_feat(186), I6 =>  inp_feat(132), I7 =>  inp_feat(36)); 
C_62_S_3_L_7_inst : LUT8 generic map(INIT => "1101110100001101110011010101011111111100010001011101111011110111110000000100000011011000110100011111000000000100111110110101111111011100110011000100000000000100010001000001000001000000000001001100000011000000010100000100010001000000110101000100000001011101") port map( O =>C_62_S_3_L_7_out, I0 =>  inp_feat(100), I1 =>  inp_feat(128), I2 =>  inp_feat(291), I3 =>  inp_feat(187), I4 =>  inp_feat(387), I5 =>  inp_feat(186), I6 =>  inp_feat(132), I7 =>  inp_feat(36)); 
C_62_S_4_L_0_inst : LUT8 generic map(INIT => "1111100110101010111100110011001111001010101110000111101100010001101010000000100010110001001100111100000100001000101100110011001100011110000000101011001010110001101100110000001111110111000000111101101110110001011101110011001111101111001000101011001100110011") port map( O =>C_62_S_4_L_0_out, I0 =>  inp_feat(60), I1 =>  inp_feat(137), I2 =>  inp_feat(130), I3 =>  inp_feat(114), I4 =>  inp_feat(398), I5 =>  inp_feat(291), I6 =>  inp_feat(69), I7 =>  inp_feat(318)); 
C_62_S_4_L_1_inst : LUT8 generic map(INIT => "0111111000111111111111111111111101011101101011010001110011111111111110001110110110111100111111110100000010000000000000001111000000010000100110111100001000110111010101010000000001000010000100010000000010011001110101110111110100000000000000000000000000000000") port map( O =>C_62_S_4_L_1_out, I0 =>  inp_feat(190), I1 =>  inp_feat(221), I2 =>  inp_feat(469), I3 =>  inp_feat(457), I4 =>  inp_feat(37), I5 =>  inp_feat(114), I6 =>  inp_feat(431), I7 =>  inp_feat(222)); 
C_62_S_4_L_2_inst : LUT8 generic map(INIT => "1100111011111110110010000100111011101110101010001100110011001110110011101010101010000100000010001100111011101110110011000100110111100000100000000000010000000000101000000100000001000000000000011101010011111000010000000000000011000000011000100000010000000000") port map( O =>C_62_S_4_L_2_out, I0 =>  inp_feat(329), I1 =>  inp_feat(483), I2 =>  inp_feat(83), I3 =>  inp_feat(472), I4 =>  inp_feat(251), I5 =>  inp_feat(398), I6 =>  inp_feat(201), I7 =>  inp_feat(256)); 
C_62_S_4_L_3_inst : LUT8 generic map(INIT => "1111111010100000101010101110111010100000101000001000000010000000001000100000000010101010000000001010000000100000100000001000000011101110111000001110111110111000101000001010000010000000000000000000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_62_S_4_L_3_out, I0 =>  inp_feat(488), I1 =>  inp_feat(172), I2 =>  inp_feat(380), I3 =>  inp_feat(396), I4 =>  inp_feat(307), I5 =>  inp_feat(209), I6 =>  inp_feat(238), I7 =>  inp_feat(472)); 
C_62_S_4_L_4_inst : LUT8 generic map(INIT => "1111101001010010000010100000000011111010001100111111000010010000010011101110001011001110000000001010110000100000110001000101001010110010101000001011001010010000111110101111101011111010111110011010101011000000100010100000000011111010111110111111101011111110") port map( O =>C_62_S_4_L_4_out, I0 =>  inp_feat(94), I1 =>  inp_feat(23), I2 =>  inp_feat(172), I3 =>  inp_feat(472), I4 =>  inp_feat(222), I5 =>  inp_feat(37), I6 =>  inp_feat(130), I7 =>  inp_feat(61)); 
C_62_S_4_L_5_inst : LUT8 generic map(INIT => "0101100111100100000000000000000011001101110011001101110100000000100101001100001001000000010000001111000101000011001000001100110011110101111111011101110111000111111111111111110101011101111111011111110011111110100001000100000001110101011101111101110111111101") port map( O =>C_62_S_4_L_5_out, I0 =>  inp_feat(408), I1 =>  inp_feat(32), I2 =>  inp_feat(342), I3 =>  inp_feat(291), I4 =>  inp_feat(182), I5 =>  inp_feat(37), I6 =>  inp_feat(336), I7 =>  inp_feat(457)); 
C_62_S_4_L_6_inst : LUT8 generic map(INIT => "1011101011011001111100101011000011111011101011111000001010100000001011110000110000100000000000000010111110100000101010110000000011011101101100011011000001000000111111110011001100110001000100000100010001000100000010000000000001010101110101010011001100000000") port map( O =>C_62_S_4_L_6_out, I0 =>  inp_feat(222), I1 =>  inp_feat(408), I2 =>  inp_feat(221), I3 =>  inp_feat(132), I4 =>  inp_feat(483), I5 =>  inp_feat(307), I6 =>  inp_feat(256), I7 =>  inp_feat(207)); 
C_62_S_4_L_7_inst : LUT8 generic map(INIT => "1100110011001110110010001100100011101110100111001110101001001001111010101110000011101010100000001011101011010000101010101000000011001000100010001100110000001000110011001100101011001000010010001100000011000000110010001000000011000100100000001110011010000000") port map( O =>C_62_S_4_L_7_out, I0 =>  inp_feat(380), I1 =>  inp_feat(238), I2 =>  inp_feat(489), I3 =>  inp_feat(336), I4 =>  inp_feat(229), I5 =>  inp_feat(291), I6 =>  inp_feat(469), I7 =>  inp_feat(196)); 
C_63_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000010000000000010000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000001000100000001000100010111000000000000000000000001000000001100000000000000010100000000000000000000000000000000000000000000") port map( O =>C_63_S_0_L_0_out, I0 =>  inp_feat(483), I1 =>  inp_feat(218), I2 =>  inp_feat(79), I3 =>  inp_feat(3), I4 =>  inp_feat(152), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_63_S_0_L_1_inst : LUT8 generic map(INIT => "0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000011001100010111000000000001010000010011000000110000000000000000000000000000000100000000000000000000001100000011000000000000000000") port map( O =>C_63_S_0_L_1_out, I0 =>  inp_feat(152), I1 =>  inp_feat(190), I2 =>  inp_feat(444), I3 =>  inp_feat(251), I4 =>  inp_feat(436), I5 =>  inp_feat(335), I6 =>  inp_feat(5), I7 =>  inp_feat(483)); 
C_63_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110010000000000000000000000000001000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_0_L_2_out, I0 =>  inp_feat(307), I1 =>  inp_feat(483), I2 =>  inp_feat(137), I3 =>  inp_feat(143), I4 =>  inp_feat(277), I5 =>  inp_feat(207), I6 =>  inp_feat(304), I7 =>  inp_feat(329)); 
C_63_S_0_L_3_inst : LUT8 generic map(INIT => "0000001100000000000000000000000000011010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010100010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_0_L_3_out, I0 =>  inp_feat(87), I1 =>  inp_feat(483), I2 =>  inp_feat(418), I3 =>  inp_feat(342), I4 =>  inp_feat(265), I5 =>  inp_feat(114), I6 =>  inp_feat(249), I7 =>  inp_feat(238)); 
C_63_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000010000000000000000000000000000000110011000000000000000000000000000000000000000000000000000000000011011100000000000000000000000000100010000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_0_L_4_out, I0 =>  inp_feat(91), I1 =>  inp_feat(36), I2 =>  inp_feat(201), I3 =>  inp_feat(408), I4 =>  inp_feat(61), I5 =>  inp_feat(23), I6 =>  inp_feat(375), I7 =>  inp_feat(152)); 
C_63_S_0_L_5_inst : LUT8 generic map(INIT => "0010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011100000111101000000100000001000000000000000010000000000000000000000000010000000000000001000110000000000000000000000000000000000") port map( O =>C_63_S_0_L_5_out, I0 =>  inp_feat(478), I1 =>  inp_feat(476), I2 =>  inp_feat(79), I3 =>  inp_feat(218), I4 =>  inp_feat(265), I5 =>  inp_feat(190), I6 =>  inp_feat(57), I7 =>  inp_feat(488)); 
C_63_S_0_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000110001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001011001000110000000000000010001100110011001100000010000000100000000000000000000000000000000000000000000000100000000000000000") port map( O =>C_63_S_0_L_6_out, I0 =>  inp_feat(201), I1 =>  inp_feat(329), I2 =>  inp_feat(467), I3 =>  inp_feat(152), I4 =>  inp_feat(322), I5 =>  inp_feat(251), I6 =>  inp_feat(190), I7 =>  inp_feat(483)); 
C_63_S_0_L_7_inst : LUT8 generic map(INIT => "0000000000000000010000001000000000000000100000001110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001000000011000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_0_L_7_out, I0 =>  inp_feat(445), I1 =>  inp_feat(190), I2 =>  inp_feat(324), I3 =>  inp_feat(437), I4 =>  inp_feat(483), I5 =>  inp_feat(226), I6 =>  inp_feat(408), I7 =>  inp_feat(91)); 
C_63_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000010000000000010000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000001000100000001000100010111000000000000000000000001000000001100000000000000010100000000000000000000000000000000000000000000") port map( O =>C_63_S_1_L_0_out, I0 =>  inp_feat(483), I1 =>  inp_feat(218), I2 =>  inp_feat(79), I3 =>  inp_feat(3), I4 =>  inp_feat(152), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_63_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000100010110000000010001000000000000000101000000000000000000000000000000111000000000000001000000010000000100000001000000000000000000000101000010110") port map( O =>C_63_S_1_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(152), I2 =>  inp_feat(483), I3 =>  inp_feat(245), I4 =>  inp_feat(488), I5 =>  inp_feat(29), I6 =>  inp_feat(187), I7 =>  inp_feat(467)); 
C_63_S_1_L_2_inst : LUT8 generic map(INIT => "0000000000000000001000000000000000000000000000000000000000000000101100110000010000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_1_L_2_out, I0 =>  inp_feat(94), I1 =>  inp_feat(483), I2 =>  inp_feat(152), I3 =>  inp_feat(100), I4 =>  inp_feat(156), I5 =>  inp_feat(190), I6 =>  inp_feat(329), I7 =>  inp_feat(288)); 
C_63_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000001000000000000000110000000000000010000000000000001100000000000000010000000000000000000000000001000100000000000000010100001000000010000000100010001000000000000000100010000000000010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_1_L_3_out, I0 =>  inp_feat(79), I1 =>  inp_feat(190), I2 =>  inp_feat(483), I3 =>  inp_feat(488), I4 =>  inp_feat(226), I5 =>  inp_feat(308), I6 =>  inp_feat(269), I7 =>  inp_feat(375)); 
C_63_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000001010000000000110101000000000000000100000100000000000000000000000000000000000000000000000000000000010000000000010000000000000000000100000000000101010000000000100111110000110000000000000000000000000000000000000000000000000") port map( O =>C_63_S_1_L_4_out, I0 =>  inp_feat(291), I1 =>  inp_feat(226), I2 =>  inp_feat(488), I3 =>  inp_feat(269), I4 =>  inp_feat(375), I5 =>  inp_feat(437), I6 =>  inp_feat(297), I7 =>  inp_feat(152)); 
C_63_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000001000000000000000000010001000100000001000100000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000000001000100010000000001110101000000000000000000000000000000000") port map( O =>C_63_S_1_L_5_out, I0 =>  inp_feat(57), I1 =>  inp_feat(272), I2 =>  inp_feat(201), I3 =>  inp_feat(283), I4 =>  inp_feat(142), I5 =>  inp_feat(424), I6 =>  inp_feat(483), I7 =>  inp_feat(128)); 
C_63_S_1_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000100000000000001101000001001000111100010000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000001000000000011010100000011000101010100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_1_L_6_out, I0 =>  inp_feat(187), I1 =>  inp_feat(201), I2 =>  inp_feat(375), I3 =>  inp_feat(170), I4 =>  inp_feat(222), I5 =>  inp_feat(483), I6 =>  inp_feat(408), I7 =>  inp_feat(416)); 
C_63_S_1_L_7_inst : LUT8 generic map(INIT => "0100000001000000010000000001000000000000000000000000000000010000000000000000000011000000010100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010100000000000001010000000100000111000000000000000000000001000000010000") port map( O =>C_63_S_1_L_7_out, I0 =>  inp_feat(483), I1 =>  inp_feat(218), I2 =>  inp_feat(408), I3 =>  inp_feat(152), I4 =>  inp_feat(488), I5 =>  inp_feat(32), I6 =>  inp_feat(182), I7 =>  inp_feat(465)); 
C_63_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000010000000000010000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000001000100000001000100010111000000000000000000000001000000001100000000000000010100000000000000000000000000000000000000000000") port map( O =>C_63_S_2_L_0_out, I0 =>  inp_feat(483), I1 =>  inp_feat(218), I2 =>  inp_feat(79), I3 =>  inp_feat(3), I4 =>  inp_feat(152), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_63_S_2_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000110100000000000011000000000000000101000000000000000000000000000001010000000000000001000000010000000100000001000000000000000000000101000001110000") port map( O =>C_63_S_2_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(152), I2 =>  inp_feat(190), I3 =>  inp_feat(496), I4 =>  inp_feat(488), I5 =>  inp_feat(29), I6 =>  inp_feat(187), I7 =>  inp_feat(467)); 
C_63_S_2_L_2_inst : LUT8 generic map(INIT => "0100000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_2_L_2_out, I0 =>  inp_feat(488), I1 =>  inp_feat(123), I2 =>  inp_feat(408), I3 =>  inp_feat(384), I4 =>  inp_feat(457), I5 =>  inp_feat(505), I6 =>  inp_feat(329), I7 =>  inp_feat(288)); 
C_63_S_2_L_3_inst : LUT8 generic map(INIT => "0000000010000110000000000100000000000000000010000000000000000000000000000100110100000000000010000000010000000100000000000000000001010010110111110000000000000000000000000000110000000000000000000000000000001000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_2_L_3_out, I0 =>  inp_feat(416), I1 =>  inp_feat(201), I2 =>  inp_feat(308), I3 =>  inp_feat(483), I4 =>  inp_feat(190), I5 =>  inp_feat(130), I6 =>  inp_feat(23), I7 =>  inp_feat(375)); 
C_63_S_2_L_4_inst : LUT8 generic map(INIT => "0001010100000000000001000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000001000111001010100100011000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_2_L_4_out, I0 =>  inp_feat(476), I1 =>  inp_feat(222), I2 =>  inp_feat(483), I3 =>  inp_feat(60), I4 =>  inp_feat(91), I5 =>  inp_feat(307), I6 =>  inp_feat(190), I7 =>  inp_feat(488)); 
C_63_S_2_L_5_inst : LUT8 generic map(INIT => "0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010111100100010000000000000010000001110000110000000000000000000000100000000000000000000000000000001000000001100000000000000000000") port map( O =>C_63_S_2_L_5_out, I0 =>  inp_feat(23), I1 =>  inp_feat(94), I2 =>  inp_feat(476), I3 =>  inp_feat(478), I4 =>  inp_feat(190), I5 =>  inp_feat(172), I6 =>  inp_feat(322), I7 =>  inp_feat(488)); 
C_63_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000100000000000001010000000000000001000000000000000100000000000000000000000000000101000000010000000000000000000000010000000000000000000000000000000100000001000001010001000100011001100000000000000000000000000000010000000100000") port map( O =>C_63_S_2_L_6_out, I0 =>  inp_feat(190), I1 =>  inp_feat(483), I2 =>  inp_feat(436), I3 =>  inp_feat(304), I4 =>  inp_feat(226), I5 =>  inp_feat(441), I6 =>  inp_feat(128), I7 =>  inp_feat(152)); 
C_63_S_2_L_7_inst : LUT8 generic map(INIT => "0000000010000000000000001000000000000000100000001000100010000000000000000000000000000000000000000000000010000000100010001000000000000000100000000000000010100000000000000000000010000000100000000000000000000000000000000000000000000000000000001110001000000000") port map( O =>C_63_S_2_L_7_out, I0 =>  inp_feat(190), I1 =>  inp_feat(387), I2 =>  inp_feat(291), I3 =>  inp_feat(335), I4 =>  inp_feat(283), I5 =>  inp_feat(483), I6 =>  inp_feat(469), I7 =>  inp_feat(294)); 
C_63_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000010000000000010000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000001000100000001000100010111000000000000000000000001000000001100000000000000010100000000000000000000000000000000000000000000") port map( O =>C_63_S_3_L_0_out, I0 =>  inp_feat(483), I1 =>  inp_feat(218), I2 =>  inp_feat(79), I3 =>  inp_feat(3), I4 =>  inp_feat(152), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_63_S_3_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000110100000000000011000000000000000101000000000000000000000000000001010000000000000001000000010000000100000001000000000000000000000101000001110000") port map( O =>C_63_S_3_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(152), I2 =>  inp_feat(190), I3 =>  inp_feat(496), I4 =>  inp_feat(488), I5 =>  inp_feat(29), I6 =>  inp_feat(187), I7 =>  inp_feat(467)); 
C_63_S_3_L_2_inst : LUT8 generic map(INIT => "0111011100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_3_L_2_out, I0 =>  inp_feat(483), I1 =>  inp_feat(437), I2 =>  inp_feat(488), I3 =>  inp_feat(49), I4 =>  inp_feat(457), I5 =>  inp_feat(388), I6 =>  inp_feat(505), I7 =>  inp_feat(288)); 
C_63_S_3_L_3_inst : LUT8 generic map(INIT => "0000001000000001000000100000001000000000000000100000000000000000000000100000001000000000001000100000001000000000000000000000000001010111000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_3_L_3_out, I0 =>  inp_feat(201), I1 =>  inp_feat(283), I2 =>  inp_feat(483), I3 =>  inp_feat(445), I4 =>  inp_feat(130), I5 =>  inp_feat(190), I6 =>  inp_feat(23), I7 =>  inp_feat(375)); 
C_63_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000001000110101000000000000000100000000000000000010000100000000000010100000000000000010000000000000000000000000000000000000000000001010000000000000001000000000000000000000000000000000000000000000") port map( O =>C_63_S_3_L_4_out, I0 =>  inp_feat(79), I1 =>  inp_feat(483), I2 =>  inp_feat(32), I3 =>  inp_feat(322), I4 =>  inp_feat(304), I5 =>  inp_feat(436), I6 =>  inp_feat(416), I7 =>  inp_feat(441)); 
C_63_S_3_L_5_inst : LUT8 generic map(INIT => "0100000011000001110100000101000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000101000001010001000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000") port map( O =>C_63_S_3_L_5_out, I0 =>  inp_feat(488), I1 =>  inp_feat(218), I2 =>  inp_feat(433), I3 =>  inp_feat(238), I4 =>  inp_feat(187), I5 =>  inp_feat(190), I6 =>  inp_feat(57), I7 =>  inp_feat(29)); 
C_63_S_3_L_6_inst : LUT8 generic map(INIT => "0000000000000000110000000100000011000000000000000101000000000000010000000000000001010100011000000000000000000000110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_3_L_6_out, I0 =>  inp_feat(488), I1 =>  inp_feat(304), I2 =>  inp_feat(207), I3 =>  inp_feat(436), I4 =>  inp_feat(483), I5 =>  inp_feat(441), I6 =>  inp_feat(152), I7 =>  inp_feat(493)); 
C_63_S_3_L_7_inst : LUT8 generic map(INIT => "0000000000000000001100000000000000110000000000000111000001000000010000000000000010000000000000000100000001000000000000000000000000110000100100000111000010000000001100000000000000110000000000000100000011000000000000000100000000000000000000000000000001000000") port map( O =>C_63_S_3_L_7_out, I0 =>  inp_feat(152), I1 =>  inp_feat(476), I2 =>  inp_feat(408), I3 =>  inp_feat(478), I4 =>  inp_feat(251), I5 =>  inp_feat(221), I6 =>  inp_feat(32), I7 =>  inp_feat(308)); 
C_63_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000010000000000010000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000001000100000001000100010111000000000000000000000001000000001100000000000000010100000000000000000000000000000000000000000000") port map( O =>C_63_S_4_L_0_out, I0 =>  inp_feat(483), I1 =>  inp_feat(218), I2 =>  inp_feat(79), I3 =>  inp_feat(3), I4 =>  inp_feat(152), I5 =>  inp_feat(190), I6 =>  inp_feat(437), I7 =>  inp_feat(488)); 
C_63_S_4_L_1_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000100000000000000000001000100000000000000000000000000010001000100010000000000000000000100000000000000010001110110011001000100010001000") port map( O =>C_63_S_4_L_1_out, I0 =>  inp_feat(396), I1 =>  inp_feat(190), I2 =>  inp_feat(475), I3 =>  inp_feat(172), I4 =>  inp_feat(437), I5 =>  inp_feat(488), I6 =>  inp_feat(187), I7 =>  inp_feat(467)); 
C_63_S_4_L_2_inst : LUT8 generic map(INIT => "0000000000000000000000000000100000001100010000001000110000001100000000000000000000000000000000000100010000010000000001000000010000000000000000000000000000001000010000000000000000000100000011000000000001000000000000000000000000001100110001010000000000000000") port map( O =>C_63_S_4_L_2_out, I0 =>  inp_feat(152), I1 =>  inp_feat(190), I2 =>  inp_feat(226), I3 =>  inp_feat(251), I4 =>  inp_feat(375), I5 =>  inp_feat(483), I6 =>  inp_feat(218), I7 =>  inp_feat(83)); 
C_63_S_4_L_3_inst : LUT8 generic map(INIT => "0001000001110000011100000011000000000000000100000000000000110010000100000000000001010000000100000000000000010000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_4_L_3_out, I0 =>  inp_feat(226), I1 =>  inp_feat(483), I2 =>  inp_feat(100), I3 =>  inp_feat(142), I4 =>  inp_feat(416), I5 =>  inp_feat(218), I6 =>  inp_feat(83), I7 =>  inp_feat(296)); 
C_63_S_4_L_4_inst : LUT8 generic map(INIT => "0000000011000000000001000000000000000000000000000101100000000000010000001100010000000000000000000100000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_4_L_4_out, I0 =>  inp_feat(483), I1 =>  inp_feat(436), I2 =>  inp_feat(130), I3 =>  inp_feat(335), I4 =>  inp_feat(79), I5 =>  inp_feat(152), I6 =>  inp_feat(418), I7 =>  inp_feat(501)); 
C_63_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010001000000001111001100000000000101010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000") port map( O =>C_63_S_4_L_5_out, I0 =>  inp_feat(187), I1 =>  inp_feat(152), I2 =>  inp_feat(218), I3 =>  inp_feat(325), I4 =>  inp_feat(38), I5 =>  inp_feat(87), I6 =>  inp_feat(190), I7 =>  inp_feat(329)); 
C_63_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000100000000000000000000000000000000000000100000000000000000000000100000000000000010000000000000000000000000000000000001001111000011110000000000000000000000000000010000000000000000100000001000100110000000000000000000001000000010000000000000000000") port map( O =>C_63_S_4_L_6_out, I0 =>  inp_feat(75), I1 =>  inp_feat(308), I2 =>  inp_feat(483), I3 =>  inp_feat(152), I4 =>  inp_feat(342), I5 =>  inp_feat(489), I6 =>  inp_feat(473), I7 =>  inp_feat(488)); 
C_63_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000001000000100000000000000000001010100000000000000000000000100010001100000000010000100000000010001000000000000000000000000000000000000000000000000000000000001000100000000000000010000000000000000000000000000000000000000000") port map( O =>C_63_S_4_L_7_out, I0 =>  inp_feat(242), I1 =>  inp_feat(79), I2 =>  inp_feat(152), I3 =>  inp_feat(342), I4 =>  inp_feat(489), I5 =>  inp_feat(473), I6 =>  inp_feat(488), I7 =>  inp_feat(442)); 
C_64_S_0_L_0_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_1_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_2_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_3_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_4_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_5_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_6_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_0_L_7_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_0_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_1_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_2_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_3_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_4_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_5_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_6_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_1_L_7_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_1_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_0_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_1_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_2_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_3_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_4_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_5_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_6_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_2_L_7_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_2_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_0_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_1_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_2_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_3_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_4_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_5_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_6_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_3_L_7_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_3_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_0_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_1_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_2_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_3_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_4_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_5_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_6_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_6_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_64_S_4_L_7_inst : LUT8 generic map(INIT => "0000000100000000000000000000000000000010101000000000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000000000000000010100010101000100000000000000000") port map( O =>C_64_S_4_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(386), I2 =>  inp_feat(14), I3 =>  inp_feat(191), I4 =>  inp_feat(302), I5 =>  inp_feat(205), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_65_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000100100000000000000100000000000000000000000100000000000000000000010100000000000000010000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101100000000000000100000000000001010000000000000") port map( O =>C_65_S_0_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_65_S_0_L_1_inst : LUT8 generic map(INIT => "0001000000010100000000011001110100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001010010010001000100001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_0_L_1_out, I0 =>  inp_feat(442), I1 =>  inp_feat(370), I2 =>  inp_feat(44), I3 =>  inp_feat(347), I4 =>  inp_feat(117), I5 =>  inp_feat(336), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_65_S_0_L_2_inst : LUT8 generic map(INIT => "0000000011000000000000000100000000000000000000000000000000000000100000000100000000000000010000000000000000000000000000000000000001000000010000001000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000") port map( O =>C_65_S_0_L_2_out, I0 =>  inp_feat(442), I1 =>  inp_feat(302), I2 =>  inp_feat(1), I3 =>  inp_feat(393), I4 =>  inp_feat(43), I5 =>  inp_feat(121), I6 =>  inp_feat(94), I7 =>  inp_feat(111)); 
C_65_S_0_L_3_inst : LUT8 generic map(INIT => "1000000010001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_0_L_3_out, I0 =>  inp_feat(388), I1 =>  inp_feat(285), I2 =>  inp_feat(105), I3 =>  inp_feat(293), I4 =>  inp_feat(283), I5 =>  inp_feat(145), I6 =>  inp_feat(172), I7 =>  inp_feat(478)); 
C_65_S_0_L_4_inst : LUT8 generic map(INIT => "0000000000000000100000000000000000000000000000000000000000000000101000000000000000000000000000000010000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_0_L_4_out, I0 =>  inp_feat(336), I1 =>  inp_feat(79), I2 =>  inp_feat(82), I3 =>  inp_feat(145), I4 =>  inp_feat(277), I5 =>  inp_feat(478), I6 =>  inp_feat(474), I7 =>  inp_feat(487)); 
C_65_S_0_L_5_inst : LUT8 generic map(INIT => "0000100000000000000000000000000000001000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000001000000010000000000000000000100010000000000000000000000000001000100000000000000000000000000000001000000000000000000000000000") port map( O =>C_65_S_0_L_5_out, I0 =>  inp_feat(179), I1 =>  inp_feat(108), I2 =>  inp_feat(168), I3 =>  inp_feat(336), I4 =>  inp_feat(89), I5 =>  inp_feat(400), I6 =>  inp_feat(303), I7 =>  inp_feat(44)); 
C_65_S_0_L_6_inst : LUT8 generic map(INIT => "0000000011000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000100000001100000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_0_L_6_out, I0 =>  inp_feat(228), I1 =>  inp_feat(154), I2 =>  inp_feat(139), I3 =>  inp_feat(241), I4 =>  inp_feat(135), I5 =>  inp_feat(168), I6 =>  inp_feat(120), I7 =>  inp_feat(442)); 
C_65_S_0_L_7_inst : LUT8 generic map(INIT => "1000001000000000101000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000001110000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_0_L_7_out, I0 =>  inp_feat(108), I1 =>  inp_feat(275), I2 =>  inp_feat(494), I3 =>  inp_feat(265), I4 =>  inp_feat(442), I5 =>  inp_feat(1), I6 =>  inp_feat(220), I7 =>  inp_feat(393)); 
C_65_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000100100000000000000100000000000000000000000100000000000000000000010100000000000000010000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101100000000000000100000000000001010000000000000") port map( O =>C_65_S_1_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_65_S_1_L_1_inst : LUT8 generic map(INIT => "0001000000100000000100000001000000000000100000001000000000110000000000000000000000000000000000000000000000000000000000000000000001000000011000000000000010110000000000000000000010010000001100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_1_L_1_out, I0 =>  inp_feat(297), I1 =>  inp_feat(442), I2 =>  inp_feat(478), I3 =>  inp_feat(474), I4 =>  inp_feat(83), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_65_S_1_L_2_inst : LUT8 generic map(INIT => "0011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_1_L_2_out, I0 =>  inp_feat(440), I1 =>  inp_feat(437), I2 =>  inp_feat(442), I3 =>  inp_feat(388), I4 =>  inp_feat(302), I5 =>  inp_feat(105), I6 =>  inp_feat(415), I7 =>  inp_feat(295)); 
C_65_S_1_L_3_inst : LUT8 generic map(INIT => "1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_1_L_3_out, I0 =>  inp_feat(193), I1 =>  inp_feat(130), I2 =>  inp_feat(448), I3 =>  inp_feat(302), I4 =>  inp_feat(9), I5 =>  inp_feat(89), I6 =>  inp_feat(462), I7 =>  inp_feat(149)); 
C_65_S_1_L_4_inst : LUT8 generic map(INIT => "1100000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_1_L_4_out, I0 =>  inp_feat(11), I1 =>  inp_feat(26), I2 =>  inp_feat(316), I3 =>  inp_feat(211), I4 =>  inp_feat(185), I5 =>  inp_feat(462), I6 =>  inp_feat(504), I7 =>  inp_feat(359)); 
C_65_S_1_L_5_inst : LUT8 generic map(INIT => "1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_1_L_5_out, I0 =>  inp_feat(40), I1 =>  inp_feat(329), I2 =>  inp_feat(462), I3 =>  inp_feat(71), I4 =>  inp_feat(130), I5 =>  inp_feat(359), I6 =>  inp_feat(139), I7 =>  inp_feat(312)); 
C_65_S_1_L_6_inst : LUT8 generic map(INIT => "0010010000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000001010110000000000000000000000000101000000000000000000000000000000000001100000000000000000000000000100010000000000000000000000000") port map( O =>C_65_S_1_L_6_out, I0 =>  inp_feat(376), I1 =>  inp_feat(442), I2 =>  inp_feat(14), I3 =>  inp_feat(89), I4 =>  inp_feat(462), I5 =>  inp_feat(132), I6 =>  inp_feat(459), I7 =>  inp_feat(468)); 
C_65_S_1_L_7_inst : LUT8 generic map(INIT => "0000000000000001000011000000000000000000000000000000000000000000011111000010000000000000000000000000000000000000000000000000000010000011000000000000000100000000000000000000000000000000000000000101110100000000010111010000000000000000000000000000000000000000") port map( O =>C_65_S_1_L_7_out, I0 =>  inp_feat(231), I1 =>  inp_feat(190), I2 =>  inp_feat(303), I3 =>  inp_feat(461), I4 =>  inp_feat(434), I5 =>  inp_feat(302), I6 =>  inp_feat(442), I7 =>  inp_feat(168)); 
C_65_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000100100000000000000100000000000000000000000100000000000000000000010100000000000000010000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101100000000000000100000000000001010000000000000") port map( O =>C_65_S_2_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_65_S_2_L_1_inst : LUT8 generic map(INIT => "0000001001000001000000100000001000000000001000000000010001000111000000000000000000000000000000000000000000000000000000000000000010100001000000000000010001000111000000000000000000001100010001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(372), I2 =>  inp_feat(442), I3 =>  inp_feat(347), I4 =>  inp_feat(393), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_65_S_2_L_2_inst : LUT8 generic map(INIT => "0100100001001100100010000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(278), I2 =>  inp_feat(442), I3 =>  inp_feat(393), I4 =>  inp_feat(241), I5 =>  inp_feat(283), I6 =>  inp_feat(89), I7 =>  inp_feat(336)); 
C_65_S_2_L_3_inst : LUT8 generic map(INIT => "0101111000000000000000000000000000000010000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(467), I2 =>  inp_feat(442), I3 =>  inp_feat(316), I4 =>  inp_feat(59), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(145)); 
C_65_S_2_L_4_inst : LUT8 generic map(INIT => "0001000011100000000100000000000000000000000000000000000000000000001100000010000010000000000000000000000000000000000000000000000001010001000000000000000000000000000000000000000000000001000000000011000010100000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_4_out, I0 =>  inp_feat(372), I1 =>  inp_feat(442), I2 =>  inp_feat(180), I3 =>  inp_feat(312), I4 =>  inp_feat(65), I5 =>  inp_feat(478), I6 =>  inp_feat(44), I7 =>  inp_feat(195)); 
C_65_S_2_L_5_inst : LUT8 generic map(INIT => "1100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_5_out, I0 =>  inp_feat(442), I1 =>  inp_feat(221), I2 =>  inp_feat(90), I3 =>  inp_feat(295), I4 =>  inp_feat(395), I5 =>  inp_feat(130), I6 =>  inp_feat(86), I7 =>  inp_feat(195)); 
C_65_S_2_L_6_inst : LUT8 generic map(INIT => "0000001010000000001000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000010000000100010000000100010001000000000000000000000000000000000001000000010000000100000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_6_out, I0 =>  inp_feat(302), I1 =>  inp_feat(235), I2 =>  inp_feat(349), I3 =>  inp_feat(44), I4 =>  inp_feat(117), I5 =>  inp_feat(450), I6 =>  inp_feat(111), I7 =>  inp_feat(393)); 
C_65_S_2_L_7_inst : LUT8 generic map(INIT => "0000001010000000010010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011101010100000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_2_L_7_out, I0 =>  inp_feat(442), I1 =>  inp_feat(434), I2 =>  inp_feat(241), I3 =>  inp_feat(168), I4 =>  inp_feat(100), I5 =>  inp_feat(462), I6 =>  inp_feat(26), I7 =>  inp_feat(393)); 
C_65_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000100100000000000000100000000000000000000000100000000000000000000010100000000000000010000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101100000000000000100000000000001010000000000000") port map( O =>C_65_S_3_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_65_S_3_L_1_inst : LUT8 generic map(INIT => "0000001001000001000000100000001000000000001000000000010001000111000000000000000000000000000000000000000000000000000000000000000010100001000000000000010001000111000000000000000000001100010001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(372), I2 =>  inp_feat(442), I3 =>  inp_feat(347), I4 =>  inp_feat(393), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_65_S_3_L_2_inst : LUT8 generic map(INIT => "0100100001001100100010000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(278), I2 =>  inp_feat(442), I3 =>  inp_feat(393), I4 =>  inp_feat(241), I5 =>  inp_feat(283), I6 =>  inp_feat(89), I7 =>  inp_feat(336)); 
C_65_S_3_L_3_inst : LUT8 generic map(INIT => "0100110001001100000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(9), I2 =>  inp_feat(442), I3 =>  inp_feat(111), I4 =>  inp_feat(59), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(145)); 
C_65_S_3_L_4_inst : LUT8 generic map(INIT => "1101000000000000000101000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_4_out, I0 =>  inp_feat(442), I1 =>  inp_feat(398), I2 =>  inp_feat(105), I3 =>  inp_feat(9), I4 =>  inp_feat(111), I5 =>  inp_feat(34), I6 =>  inp_feat(265), I7 =>  inp_feat(195)); 
C_65_S_3_L_5_inst : LUT8 generic map(INIT => "0000100000000000000000000000000010001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_5_out, I0 =>  inp_feat(336), I1 =>  inp_feat(221), I2 =>  inp_feat(312), I3 =>  inp_feat(209), I4 =>  inp_feat(478), I5 =>  inp_feat(44), I6 =>  inp_feat(171), I7 =>  inp_feat(195)); 
C_65_S_3_L_6_inst : LUT8 generic map(INIT => "0000001000001010000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000010101010101010000100000000000000000000000000000000000000000000001010100001000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_6_out, I0 =>  inp_feat(180), I1 =>  inp_feat(434), I2 =>  inp_feat(437), I3 =>  inp_feat(14), I4 =>  inp_feat(171), I5 =>  inp_feat(463), I6 =>  inp_feat(347), I7 =>  inp_feat(442)); 
C_65_S_3_L_7_inst : LUT8 generic map(INIT => "0100000001000000000000000000000011001000000000000000000000000000010000000000000000000000000000000100001000000000000000000000000011000000000000000000000000000000100010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_3_L_7_out, I0 =>  inp_feat(241), I1 =>  inp_feat(265), I2 =>  inp_feat(108), I3 =>  inp_feat(494), I4 =>  inp_feat(7), I5 =>  inp_feat(372), I6 =>  inp_feat(505), I7 =>  inp_feat(60)); 
C_65_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000100100000000000000100000000000000000000000100000000000000000000010100000000000000010000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101100000000000000100000000000001010000000000000") port map( O =>C_65_S_4_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_65_S_4_L_1_inst : LUT8 generic map(INIT => "0000001001000001000000100000001000000000001000000000010001000111000000000000000000000000000000000000000000000000000000000000000010100001000000000000010001000111000000000000000000001100010001000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_4_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(372), I2 =>  inp_feat(442), I3 =>  inp_feat(347), I4 =>  inp_feat(393), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_65_S_4_L_2_inst : LUT8 generic map(INIT => "0100100001001100100010000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_4_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(278), I2 =>  inp_feat(442), I3 =>  inp_feat(393), I4 =>  inp_feat(241), I5 =>  inp_feat(283), I6 =>  inp_feat(89), I7 =>  inp_feat(336)); 
C_65_S_4_L_3_inst : LUT8 generic map(INIT => "0100110001001100000000000000001000000000000000000000000000001000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_4_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(139), I2 =>  inp_feat(442), I3 =>  inp_feat(293), I4 =>  inp_feat(108), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(145)); 
C_65_S_4_L_4_inst : LUT8 generic map(INIT => "1011001100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_65_S_4_L_4_out, I0 =>  inp_feat(33), I1 =>  inp_feat(442), I2 =>  inp_feat(172), I3 =>  inp_feat(478), I4 =>  inp_feat(329), I5 =>  inp_feat(390), I6 =>  inp_feat(424), I7 =>  inp_feat(34)); 
C_65_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000010000000000000001001100000000001000100000000000100000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000010001000000000011000100000000000100000000000000000000000000000001000100000000000100000000000000") port map( O =>C_65_S_4_L_5_out, I0 =>  inp_feat(499), I1 =>  inp_feat(452), I2 =>  inp_feat(434), I3 =>  inp_feat(145), I4 =>  inp_feat(14), I5 =>  inp_feat(241), I6 =>  inp_feat(112), I7 =>  inp_feat(44)); 
C_65_S_4_L_6_inst : LUT8 generic map(INIT => "0000001000000000100000000000000010000000000000000000000000000000000010100000100000000000000000000000000000000000000000000000000010001100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000100010000000000000000000000000") port map( O =>C_65_S_4_L_6_out, I0 =>  inp_feat(478), I1 =>  inp_feat(191), I2 =>  inp_feat(440), I3 =>  inp_feat(336), I4 =>  inp_feat(449), I5 =>  inp_feat(112), I6 =>  inp_feat(44), I7 =>  inp_feat(442)); 
C_65_S_4_L_7_inst : LUT8 generic map(INIT => "0000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000110000001000000000000000000000000100000000000000000000000000000010001000000000000000000000000000") port map( O =>C_65_S_4_L_7_out, I0 =>  inp_feat(331), I1 =>  inp_feat(494), I2 =>  inp_feat(180), I3 =>  inp_feat(349), I4 =>  inp_feat(7), I5 =>  inp_feat(364), I6 =>  inp_feat(372), I7 =>  inp_feat(49)); 
C_66_S_0_L_0_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_0_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_1_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_1_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_2_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_2_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_3_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_3_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_4_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_4_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_5_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_5_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_6_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_6_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_0_L_7_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_0_L_7_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_0_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_0_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_1_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_1_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_2_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_2_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_3_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_3_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_4_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_4_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_5_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_5_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_6_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_6_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_1_L_7_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_1_L_7_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_0_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_0_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_1_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_1_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_2_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_2_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_3_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_3_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_4_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_4_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_5_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_5_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_6_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_6_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_2_L_7_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_2_L_7_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_0_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_0_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_1_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_1_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_2_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_2_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_3_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_3_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_4_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_4_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_5_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_5_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_6_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_6_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_3_L_7_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_3_L_7_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_0_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_0_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_1_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_1_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_2_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_2_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_3_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_3_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_4_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_4_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_5_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_5_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_6_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_6_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_66_S_4_L_7_inst : LUT8 generic map(INIT => "0001010000000000000010010000000000000000000000000010000000000000000000000000000000100010000000000000000000000000101000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000001000100000000000101010000000001010001000000000") port map( O =>C_66_S_4_L_7_out, I0 =>  inp_feat(16), I1 =>  inp_feat(231), I2 =>  inp_feat(219), I3 =>  inp_feat(302), I4 =>  inp_feat(205), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_67_S_0_L_0_inst : LUT8 generic map(INIT => "1111001110110000111101000000000011111000010000001101100000000000011100001010000000000000000000000000000000000000000000000000000011110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_0_L_0_out, I0 =>  inp_feat(437), I1 =>  inp_feat(149), I2 =>  inp_feat(67), I3 =>  inp_feat(44), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_67_S_0_L_1_inst : LUT8 generic map(INIT => "1111001111110000000000001000000011100000101000001110010010000000101111111000000000100000000000001010000000000000011000000000000000110000000000000010000000000000000000000000000011100000000000001010000010000000101100000000000000100000000000001011000000000000") port map( O =>C_67_S_0_L_1_out, I0 =>  inp_feat(474), I1 =>  inp_feat(273), I2 =>  inp_feat(231), I3 =>  inp_feat(330), I4 =>  inp_feat(11), I5 =>  inp_feat(4), I6 =>  inp_feat(46), I7 =>  inp_feat(312)); 
C_67_S_0_L_2_inst : LUT8 generic map(INIT => "0110111011101010100010101110101010101000101010001000100000000000011011001110101011101010110010101010000000100000000010000000000011111000111111101010101000000010100010001010100010001000000000000111000000000000100000000000000000100000000000000000000000000000") port map( O =>C_67_S_0_L_2_out, I0 =>  inp_feat(17), I1 =>  inp_feat(26), I2 =>  inp_feat(336), I3 =>  inp_feat(478), I4 =>  inp_feat(371), I5 =>  inp_feat(141), I6 =>  inp_feat(388), I7 =>  inp_feat(221)); 
C_67_S_0_L_3_inst : LUT8 generic map(INIT => "0110100011101000111011101010000011101110010001000010101010100000101010101010100011101110100010101010101000000000001000100000000011000000101010001010110010100000000000000000000000100000001000001111100010111000111011101010101000000000000000000000000000000000") port map( O =>C_67_S_0_L_3_out, I0 =>  inp_feat(192), I1 =>  inp_feat(211), I2 =>  inp_feat(149), I3 =>  inp_feat(171), I4 =>  inp_feat(26), I5 =>  inp_feat(395), I6 =>  inp_feat(478), I7 =>  inp_feat(365)); 
C_67_S_0_L_4_inst : LUT8 generic map(INIT => "0111101111101000101010101100100011100010110000000000001000000000111111111100100011111111110010001001000010000000000000000000000010000000101000001111101010101000100000001000000000000000100000001000000000000000000000000000000010000000100000000000000000000000") port map( O =>C_67_S_0_L_4_out, I0 =>  inp_feat(223), I1 =>  inp_feat(89), I2 =>  inp_feat(450), I3 =>  inp_feat(336), I4 =>  inp_feat(478), I5 =>  inp_feat(337), I6 =>  inp_feat(221), I7 =>  inp_feat(271)); 
C_67_S_0_L_5_inst : LUT8 generic map(INIT => "0111111100101100111110000000000011111111000000001100101000000000101100000000000011010000000000001111111100000000110000000000000010111111101011110010101000000000101110000000000010001000000000001011001000000000100000001000000010110000000000001000000010000000") port map( O =>C_67_S_0_L_5_out, I0 =>  inp_feat(130), I1 =>  inp_feat(171), I2 =>  inp_feat(82), I3 =>  inp_feat(168), I4 =>  inp_feat(145), I5 =>  inp_feat(478), I6 =>  inp_feat(387), I7 =>  inp_feat(472)); 
C_67_S_0_L_6_inst : LUT8 generic map(INIT => "1110110011001100010011000000000010101100000010000000100000000000110011001000100001000100000000001000100000000000000000000000000000001100000011000100000000000000000010000000100000000000000000001101000010001100010100000000100000000000000000000000000000000000") port map( O =>C_67_S_0_L_6_out, I0 =>  inp_feat(201), I1 =>  inp_feat(168), I2 =>  inp_feat(221), I3 =>  inp_feat(455), I4 =>  inp_feat(111), I5 =>  inp_feat(401), I6 =>  inp_feat(80), I7 =>  inp_feat(68)); 
C_67_S_0_L_7_inst : LUT8 generic map(INIT => "1111000011000000110000001100000011110000111010001010100011010000000000001100000010101000110000000000000010100000100010001000000000110000100110000000000001010000101100001101100000010000011100000000000011000000000000000000000000000000111100000000000011000000") port map( O =>C_67_S_0_L_7_out, I0 =>  inp_feat(0), I1 =>  inp_feat(7), I2 =>  inp_feat(393), I3 =>  inp_feat(180), I4 =>  inp_feat(26), I5 =>  inp_feat(478), I6 =>  inp_feat(68), I7 =>  inp_feat(474)); 
C_67_S_1_L_0_inst : LUT8 generic map(INIT => "1111001110110000111101000000000011111000010000001101100000000000011100001010000000000000000000000000000000000000000000000000000011110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_1_L_0_out, I0 =>  inp_feat(437), I1 =>  inp_feat(149), I2 =>  inp_feat(67), I3 =>  inp_feat(44), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_67_S_1_L_1_inst : LUT8 generic map(INIT => "1111001111110000000000001000000011100000101000001110010010000000101111111000000000100000000000001010000000000000011000000000000000110000000000000010000000000000000000000000000011100000000000001010000010000000101100000000000000100000000000001011000000000000") port map( O =>C_67_S_1_L_1_out, I0 =>  inp_feat(474), I1 =>  inp_feat(273), I2 =>  inp_feat(231), I3 =>  inp_feat(330), I4 =>  inp_feat(11), I5 =>  inp_feat(4), I6 =>  inp_feat(46), I7 =>  inp_feat(312)); 
C_67_S_1_L_2_inst : LUT8 generic map(INIT => "0110111011101010100010101110101010101000101010001000100000000000011011001110101011101010110010101010000000100000000010000000000011111000111111101010101000000010100010001010100010001000000000000111000000000000100000000000000000100000000000000000000000000000") port map( O =>C_67_S_1_L_2_out, I0 =>  inp_feat(17), I1 =>  inp_feat(26), I2 =>  inp_feat(336), I3 =>  inp_feat(478), I4 =>  inp_feat(371), I5 =>  inp_feat(141), I6 =>  inp_feat(388), I7 =>  inp_feat(221)); 
C_67_S_1_L_3_inst : LUT8 generic map(INIT => "0110100011101000111011101010000011101110010001000010101010100000101010101010100011101110100010101010101000000000001000100000000011000000101010001010110010100000000000000000000000100000001000001111100010111000111011101010101000000000000000000000000000000000") port map( O =>C_67_S_1_L_3_out, I0 =>  inp_feat(192), I1 =>  inp_feat(211), I2 =>  inp_feat(149), I3 =>  inp_feat(171), I4 =>  inp_feat(26), I5 =>  inp_feat(395), I6 =>  inp_feat(478), I7 =>  inp_feat(365)); 
C_67_S_1_L_4_inst : LUT8 generic map(INIT => "0111101111101000101010101100100011100010110000000000001000000000111111111100100011111111110010001001000010000000000000000000000010000000101000001111101010101000100000001000000000000000100000001000000000000000000000000000000010000000100000000000000000000000") port map( O =>C_67_S_1_L_4_out, I0 =>  inp_feat(223), I1 =>  inp_feat(89), I2 =>  inp_feat(450), I3 =>  inp_feat(336), I4 =>  inp_feat(478), I5 =>  inp_feat(337), I6 =>  inp_feat(221), I7 =>  inp_feat(271)); 
C_67_S_1_L_5_inst : LUT8 generic map(INIT => "0111111100101100111110000000000011111111000000001100101000000000101100000000000011010000000000001111111100000000110000000000000010111111101011110010101000000000101110000000000010001000000000001011001000000000100000001000000010110000000000001000000010000000") port map( O =>C_67_S_1_L_5_out, I0 =>  inp_feat(130), I1 =>  inp_feat(171), I2 =>  inp_feat(82), I3 =>  inp_feat(168), I4 =>  inp_feat(145), I5 =>  inp_feat(478), I6 =>  inp_feat(387), I7 =>  inp_feat(472)); 
C_67_S_1_L_6_inst : LUT8 generic map(INIT => "1111111111011111010011011100110011001110010010000100110011000000110111100000000000000100110000001100000001000000110011001100000000001000000010000000000000000000000010000000100000000000000000001100111000000000110011010000000000000000000000000000000000000000") port map( O =>C_67_S_1_L_6_out, I0 =>  inp_feat(478), I1 =>  inp_feat(117), I2 =>  inp_feat(221), I3 =>  inp_feat(325), I4 =>  inp_feat(474), I5 =>  inp_feat(401), I6 =>  inp_feat(80), I7 =>  inp_feat(68)); 
C_67_S_1_L_7_inst : LUT8 generic map(INIT => "1111111111111110000101001111111011111111111111000000000000110100111101111010101000001100110011001111111100000000000000000000010010000000100010000000000000000000100011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_1_L_7_out, I0 =>  inp_feat(469), I1 =>  inp_feat(180), I2 =>  inp_feat(303), I3 =>  inp_feat(478), I4 =>  inp_feat(386), I5 =>  inp_feat(21), I6 =>  inp_feat(312), I7 =>  inp_feat(168)); 
C_67_S_2_L_0_inst : LUT8 generic map(INIT => "1111001110110000111101000000000011111000010000001101100000000000011100001010000000000000000000000000000000000000000000000000000011110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_2_L_0_out, I0 =>  inp_feat(437), I1 =>  inp_feat(149), I2 =>  inp_feat(67), I3 =>  inp_feat(44), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_67_S_2_L_1_inst : LUT8 generic map(INIT => "1111001111110000000000001000000011100000101000001110010010000000101111111000000000100000000000001010000000000000011000000000000000110000000000000010000000000000000000000000000011100000000000001010000010000000101100000000000000100000000000001011000000000000") port map( O =>C_67_S_2_L_1_out, I0 =>  inp_feat(474), I1 =>  inp_feat(273), I2 =>  inp_feat(231), I3 =>  inp_feat(330), I4 =>  inp_feat(11), I5 =>  inp_feat(4), I6 =>  inp_feat(46), I7 =>  inp_feat(312)); 
C_67_S_2_L_2_inst : LUT8 generic map(INIT => "0110111011101010100010101110101010101000101010001000100000000000011011001110101011101010110010101010000000100000000010000000000011111000111111101010101000000010100010001010100010001000000000000111000000000000100000000000000000100000000000000000000000000000") port map( O =>C_67_S_2_L_2_out, I0 =>  inp_feat(17), I1 =>  inp_feat(26), I2 =>  inp_feat(336), I3 =>  inp_feat(478), I4 =>  inp_feat(371), I5 =>  inp_feat(141), I6 =>  inp_feat(388), I7 =>  inp_feat(221)); 
C_67_S_2_L_3_inst : LUT8 generic map(INIT => "0110100011101000111011101010000011101110010001000010101010100000101010101010100011101110100010101010101000000000001000100000000011000000101010001010110010100000000000000000000000100000001000001111100010111000111011101010101000000000000000000000000000000000") port map( O =>C_67_S_2_L_3_out, I0 =>  inp_feat(192), I1 =>  inp_feat(211), I2 =>  inp_feat(149), I3 =>  inp_feat(171), I4 =>  inp_feat(26), I5 =>  inp_feat(395), I6 =>  inp_feat(478), I7 =>  inp_feat(365)); 
C_67_S_2_L_4_inst : LUT8 generic map(INIT => "0111101111101000101010101100100011100010110000000000001000000000111111111100100011111111110010001001000010000000000000000000000010000000101000001111101010101000100000001000000000000000100000001000000000000000000000000000000010000000100000000000000000000000") port map( O =>C_67_S_2_L_4_out, I0 =>  inp_feat(223), I1 =>  inp_feat(89), I2 =>  inp_feat(450), I3 =>  inp_feat(336), I4 =>  inp_feat(478), I5 =>  inp_feat(337), I6 =>  inp_feat(221), I7 =>  inp_feat(271)); 
C_67_S_2_L_5_inst : LUT8 generic map(INIT => "0111111100101100111110000000000011111111000000001100101000000000101100000000000011010000000000001111111100000000110000000000000010111111101011110010101000000000101110000000000010001000000000001011001000000000100000001000000010110000000000001000000010000000") port map( O =>C_67_S_2_L_5_out, I0 =>  inp_feat(130), I1 =>  inp_feat(171), I2 =>  inp_feat(82), I3 =>  inp_feat(168), I4 =>  inp_feat(145), I5 =>  inp_feat(478), I6 =>  inp_feat(387), I7 =>  inp_feat(472)); 
C_67_S_2_L_6_inst : LUT8 generic map(INIT => "1100110011111111110011001111011101011100101011110101110000000100110011001100110000001000000000000000100000001000000010000000000001000000100010000000000010100000000000000000000000000000000000001100010010001000000000000000000000001010000011110000000000000000") port map( O =>C_67_S_2_L_6_out, I0 =>  inp_feat(285), I1 =>  inp_feat(14), I2 =>  inp_feat(324), I3 =>  inp_feat(221), I4 =>  inp_feat(325), I5 =>  inp_feat(474), I6 =>  inp_feat(80), I7 =>  inp_feat(68)); 
C_67_S_2_L_7_inst : LUT8 generic map(INIT => "1010101011101010000010001010001010110011101110110000000000000000001010011010100000000000000010001010001110110010000000000000000000100000101000000000000000000000101000001010000000000000000000000000000000000000000000000000000010100000001000000000000000000000") port map( O =>C_67_S_2_L_7_out, I0 =>  inp_feat(454), I1 =>  inp_feat(145), I2 =>  inp_feat(223), I3 =>  inp_feat(478), I4 =>  inp_feat(112), I5 =>  inp_feat(26), I6 =>  inp_feat(93), I7 =>  inp_feat(393)); 
C_67_S_3_L_0_inst : LUT8 generic map(INIT => "1111001110110000111101000000000011111000010000001101100000000000011100001010000000000000000000000000000000000000000000000000000011110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_3_L_0_out, I0 =>  inp_feat(437), I1 =>  inp_feat(149), I2 =>  inp_feat(67), I3 =>  inp_feat(44), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_67_S_3_L_1_inst : LUT8 generic map(INIT => "1111001111110000000000001000000011100000101000001110010010000000101111111000000000100000000000001010000000000000011000000000000000110000000000000010000000000000000000000000000011100000000000001010000010000000101100000000000000100000000000001011000000000000") port map( O =>C_67_S_3_L_1_out, I0 =>  inp_feat(474), I1 =>  inp_feat(273), I2 =>  inp_feat(231), I3 =>  inp_feat(330), I4 =>  inp_feat(11), I5 =>  inp_feat(4), I6 =>  inp_feat(46), I7 =>  inp_feat(312)); 
C_67_S_3_L_2_inst : LUT8 generic map(INIT => "0110111011101010100010101110101010101000101010001000100000000000011011001110101011101010110010101010000000100000000010000000000011111000111111101010101000000010100010001010100010001000000000000111000000000000100000000000000000100000000000000000000000000000") port map( O =>C_67_S_3_L_2_out, I0 =>  inp_feat(17), I1 =>  inp_feat(26), I2 =>  inp_feat(336), I3 =>  inp_feat(478), I4 =>  inp_feat(371), I5 =>  inp_feat(141), I6 =>  inp_feat(388), I7 =>  inp_feat(221)); 
C_67_S_3_L_3_inst : LUT8 generic map(INIT => "0110100011101000111011101010000011101110010001000010101010100000101010101010100011101110100010101010101000000000001000100000000011000000101010001010110010100000000000000000000000100000001000001111100010111000111011101010101000000000000000000000000000000000") port map( O =>C_67_S_3_L_3_out, I0 =>  inp_feat(192), I1 =>  inp_feat(211), I2 =>  inp_feat(149), I3 =>  inp_feat(171), I4 =>  inp_feat(26), I5 =>  inp_feat(395), I6 =>  inp_feat(478), I7 =>  inp_feat(365)); 
C_67_S_3_L_4_inst : LUT8 generic map(INIT => "0111101111101000101010101100100011100010110000000000001000000000111111111100100011111111110010001001000010000000000000000000000010000000101000001111101010101000100000001000000000000000100000001000000000000000000000000000000010000000100000000000000000000000") port map( O =>C_67_S_3_L_4_out, I0 =>  inp_feat(223), I1 =>  inp_feat(89), I2 =>  inp_feat(450), I3 =>  inp_feat(336), I4 =>  inp_feat(478), I5 =>  inp_feat(337), I6 =>  inp_feat(221), I7 =>  inp_feat(271)); 
C_67_S_3_L_5_inst : LUT8 generic map(INIT => "0111111100101100111110000000000011111111000000001100101000000000101100000000000011010000000000001111111100000000110000000000000010111111101011110010101000000000101110000000000010001000000000001011001000000000100000001000000010110000000000001000000010000000") port map( O =>C_67_S_3_L_5_out, I0 =>  inp_feat(130), I1 =>  inp_feat(171), I2 =>  inp_feat(82), I3 =>  inp_feat(168), I4 =>  inp_feat(145), I5 =>  inp_feat(478), I6 =>  inp_feat(387), I7 =>  inp_feat(472)); 
C_67_S_3_L_6_inst : LUT8 generic map(INIT => "1011101111101011100010111110001010101010111100101010001011100010001000000100000010100010011000101010000011100010001000101110001000000010101000001000000000110010000000000010001000000000001100100010000000100000000000000000000000000010001100100000000000000010") port map( O =>C_67_S_3_L_6_out, I0 =>  inp_feat(148), I1 =>  inp_feat(4), I2 =>  inp_feat(483), I3 =>  inp_feat(351), I4 =>  inp_feat(145), I5 =>  inp_feat(478), I6 =>  inp_feat(474), I7 =>  inp_feat(68)); 
C_67_S_3_L_7_inst : LUT8 generic map(INIT => "1011101111101011100010111110001010101010111100101010001011100010001000000100000010100010011000101010000011100010001000101110001000000010101000001000000000110010000000000010001000000000001100100010000000100000000000000000000000000010001100100000000000000010") port map( O =>C_67_S_3_L_7_out, I0 =>  inp_feat(148), I1 =>  inp_feat(4), I2 =>  inp_feat(483), I3 =>  inp_feat(351), I4 =>  inp_feat(145), I5 =>  inp_feat(478), I6 =>  inp_feat(474), I7 =>  inp_feat(68)); 
C_67_S_4_L_0_inst : LUT8 generic map(INIT => "1111001110110000111101000000000011111000010000001101100000000000011100001010000000000000000000000000000000000000000000000000000011110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_4_L_0_out, I0 =>  inp_feat(437), I1 =>  inp_feat(149), I2 =>  inp_feat(67), I3 =>  inp_feat(44), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_67_S_4_L_1_inst : LUT8 generic map(INIT => "1111111011100000111011001010000000000000000000001000100000000000111110101011000010101000101000000000000000000000101010100000000000100000101000001010000010100000000000000000000000000000000000001110000011100000000000001010000000000000000000000000000000000000") port map( O =>C_67_S_4_L_1_out, I0 =>  inp_feat(440), I1 =>  inp_feat(460), I2 =>  inp_feat(111), I3 =>  inp_feat(43), I4 =>  inp_feat(328), I5 =>  inp_feat(231), I6 =>  inp_feat(46), I7 =>  inp_feat(312)); 
C_67_S_4_L_2_inst : LUT8 generic map(INIT => "1110001010101010101000101000101000000000000000001100000000000000100000001000100010000000100010000000000000000000000000000000000010100010101010101010001010001010000000000000000000000000000000001011100010101000101000001000000000000000000000000000000000000000") port map( O =>C_67_S_4_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(428), I2 =>  inp_feat(241), I3 =>  inp_feat(154), I4 =>  inp_feat(450), I5 =>  inp_feat(393), I6 =>  inp_feat(334), I7 =>  inp_feat(509)); 
C_67_S_4_L_3_inst : LUT8 generic map(INIT => "1111001110110000101110110000000011100000000000000000000000000000111000001000000000100000000000000000000000000000000000000000000011111111001100001011011100000000100010000000000000000000000000000010100000000000000000100000000000000000000000000000000000000000") port map( O =>C_67_S_4_L_3_out, I0 =>  inp_feat(123), I1 =>  inp_feat(180), I2 =>  inp_feat(43), I3 =>  inp_feat(231), I4 =>  inp_feat(205), I5 =>  inp_feat(83), I6 =>  inp_feat(117), I7 =>  inp_feat(509)); 
C_67_S_4_L_4_inst : LUT8 generic map(INIT => "0110101011001010100011001100000011101000110000001000000011000000111110001100000011001100100000001100110011001000100000001000000001111010101110100000000010000000000000001000000000000000100000001111101011101000110000001100000011101000100010001000000010000000") port map( O =>C_67_S_4_L_4_out, I0 =>  inp_feat(5), I1 =>  inp_feat(17), I2 =>  inp_feat(26), I3 =>  inp_feat(329), I4 =>  inp_feat(141), I5 =>  inp_feat(336), I6 =>  inp_feat(478), I7 =>  inp_feat(211)); 
C_67_S_4_L_5_inst : LUT8 generic map(INIT => "1101110011011100110011001101000000001100100000000000110000000000110110001100000000000000110000000100000010000000000000000000000001001100110110001100110011010000000000000000000010000000100000001100100000000000010000000000000000000000000000000000000000000000") port map( O =>C_67_S_4_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(393), I2 =>  inp_feat(444), I3 =>  inp_feat(26), I4 =>  inp_feat(120), I5 =>  inp_feat(349), I6 =>  inp_feat(225), I7 =>  inp_feat(372)); 
C_67_S_4_L_6_inst : LUT8 generic map(INIT => "1111111111011101110011111100110111000000000000001100000100000000111111110101000011000000110000000000000000000000000000000000000000001000000010001000000000000000000000000000000000000000000000001000101100000000100000000000000000000000000000000000000000000000") port map( O =>C_67_S_4_L_6_out, I0 =>  inp_feat(145), I1 =>  inp_feat(241), I2 =>  inp_feat(84), I3 =>  inp_feat(297), I4 =>  inp_feat(478), I5 =>  inp_feat(231), I6 =>  inp_feat(440), I7 =>  inp_feat(347)); 
C_67_S_4_L_7_inst : LUT8 generic map(INIT => "1110111011001100011011000000000011101010110000001000000000000000100010100000100000000000000000000000100000000000000000000000000010101000101000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_67_S_4_L_7_out, I0 =>  inp_feat(43), I1 =>  inp_feat(148), I2 =>  inp_feat(123), I3 =>  inp_feat(425), I4 =>  inp_feat(349), I5 =>  inp_feat(372), I6 =>  inp_feat(168), I7 =>  inp_feat(231)); 
C_68_S_0_L_0_inst : LUT8 generic map(INIT => "1110110110101101000010001000110011001000100010001000000010001000100000010000000100000000000000000000000000000000000000000000000010001100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_0_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_68_S_0_L_1_inst : LUT8 generic map(INIT => "1110100011000000101100000000000011110000111000000000000000000000110000001100000010000000000000001111000011000000001000000000000000000000000000000000000000000000101100000000000000000000000000001110000001000000000000000000000001110010010000000000000000000000") port map( O =>C_68_S_0_L_1_out, I0 =>  inp_feat(442), I1 =>  inp_feat(370), I2 =>  inp_feat(44), I3 =>  inp_feat(347), I4 =>  inp_feat(117), I5 =>  inp_feat(336), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_68_S_0_L_2_inst : LUT8 generic map(INIT => "1111111100001000101100000000000010101000000000001010000000000000001010000000000010100000000000001010100000001000101000000000000010111111000000000000000000000000000010000000100000000000000000000000100000000000000000000000000010001000000010000000000000000000") port map( O =>C_68_S_0_L_2_out, I0 =>  inp_feat(442), I1 =>  inp_feat(302), I2 =>  inp_feat(1), I3 =>  inp_feat(393), I4 =>  inp_feat(43), I5 =>  inp_feat(121), I6 =>  inp_feat(94), I7 =>  inp_feat(111)); 
C_68_S_0_L_3_inst : LUT8 generic map(INIT => "0111110100100111111010101000000011000000111111111000000010000000110011000000000011001110000000001110000000000000110000000000000011111010101010111010101010101000011000001111111100000000100000001100101000001010000010100000000000000001001000100000000000000000") port map( O =>C_68_S_0_L_3_out, I0 =>  inp_feat(388), I1 =>  inp_feat(285), I2 =>  inp_feat(105), I3 =>  inp_feat(293), I4 =>  inp_feat(283), I5 =>  inp_feat(145), I6 =>  inp_feat(172), I7 =>  inp_feat(478)); 
C_68_S_0_L_4_inst : LUT8 generic map(INIT => "1111110111001100000010001000100011111101110010000000100010001000010110010100000000001000110010001101110111011001110011010100100010000101101000001000000010100000101000001010000010000000101000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_68_S_0_L_4_out, I0 =>  inp_feat(336), I1 =>  inp_feat(79), I2 =>  inp_feat(82), I3 =>  inp_feat(145), I4 =>  inp_feat(277), I5 =>  inp_feat(478), I6 =>  inp_feat(474), I7 =>  inp_feat(487)); 
C_68_S_0_L_5_inst : LUT8 generic map(INIT => "1111000011111000111100100100000011100000100010001011000000000000011100001111000010100010000000001011000011110000000000000000000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_0_L_5_out, I0 =>  inp_feat(179), I1 =>  inp_feat(108), I2 =>  inp_feat(168), I3 =>  inp_feat(336), I4 =>  inp_feat(89), I5 =>  inp_feat(400), I6 =>  inp_feat(303), I7 =>  inp_feat(44)); 
C_68_S_0_L_6_inst : LUT8 generic map(INIT => "1111111100110011111011001010000001001100000000001100110000000000111100011010000110100000101000001000000000000000100000000000000000100111000001110000000000000000000001000000000000000000000000001010010100000011000000000000000000000000000000000000000000000000") port map( O =>C_68_S_0_L_6_out, I0 =>  inp_feat(228), I1 =>  inp_feat(154), I2 =>  inp_feat(139), I3 =>  inp_feat(241), I4 =>  inp_feat(135), I5 =>  inp_feat(168), I6 =>  inp_feat(120), I7 =>  inp_feat(442)); 
C_68_S_0_L_7_inst : LUT8 generic map(INIT => "0110110111101101010001010000000011001111110011011000010010000000000011111100100011001111010000001000000011000000010001000100000000000000000000000000000000000000110001010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_0_L_7_out, I0 =>  inp_feat(108), I1 =>  inp_feat(275), I2 =>  inp_feat(494), I3 =>  inp_feat(265), I4 =>  inp_feat(442), I5 =>  inp_feat(1), I6 =>  inp_feat(220), I7 =>  inp_feat(393)); 
C_68_S_1_L_0_inst : LUT8 generic map(INIT => "1110110110101101000010001000110011001000100010001000000010001000100000010000000100000000000000000000000000000000000000000000000010001100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_1_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_68_S_1_L_1_inst : LUT8 generic map(INIT => "1110111011001110110011000000010011001100000010010000000000000000111010100100111000100000000000001000000000000100000000000000000010000100000011000010000000000000000000000000000000000000000000001110110011001100001000000000000000000000000000000000000000000000") port map( O =>C_68_S_1_L_1_out, I0 =>  inp_feat(297), I1 =>  inp_feat(442), I2 =>  inp_feat(478), I3 =>  inp_feat(474), I4 =>  inp_feat(83), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_68_S_1_L_2_inst : LUT8 generic map(INIT => "1000101000001000111011100000100010101111000000001010111100000000101010000000100010101010000010001010111100000000101011110000000010101000101011101010100000101000101000000000000010100000000000001010100000001000101000000000000000000000000000000000000000000000") port map( O =>C_68_S_1_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(303), I2 =>  inp_feat(331), I3 =>  inp_feat(442), I4 =>  inp_feat(388), I5 =>  inp_feat(346), I6 =>  inp_feat(478), I7 =>  inp_feat(418)); 
C_68_S_1_L_3_inst : LUT8 generic map(INIT => "1111110101010000100000000000000001110000000100001010000010000000111100110101000011000000000000001111001101010000111000000000000010100000000000001000000000000000101000000000000011100000110000001000001100000000100000000000000010011001000000001110000011000000") port map( O =>C_68_S_1_L_3_out, I0 =>  inp_feat(462), I1 =>  inp_feat(172), I2 =>  inp_feat(264), I3 =>  inp_feat(168), I4 =>  inp_feat(58), I5 =>  inp_feat(437), I6 =>  inp_feat(344), I7 =>  inp_feat(145)); 
C_68_S_1_L_4_inst : LUT8 generic map(INIT => "1100110011011000110001001000100001000100100010001100010010001000111011001100100010100000100000000000000010001000000000001000000001001100110000000000000000000000000000000000000000000000000000001110110011001000101000001000000000001000100010000000000000000000") port map( O =>C_68_S_1_L_4_out, I0 =>  inp_feat(336), I1 =>  inp_feat(44), I2 =>  inp_feat(177), I3 =>  inp_feat(26), I4 =>  inp_feat(395), I5 =>  inp_feat(345), I6 =>  inp_feat(1), I7 =>  inp_feat(111)); 
C_68_S_1_L_5_inst : LUT8 generic map(INIT => "1110111001001000111000100000000011100100110000001100000000000000001010000000001000000000000000001111001000000000000000000000000000101111001000110010001000000000111111111111011100000000000000000000001000000000000000000000000011110010000000000000000000000000") port map( O =>C_68_S_1_L_5_out, I0 =>  inp_feat(436), I1 =>  inp_feat(278), I2 =>  inp_feat(242), I3 =>  inp_feat(132), I4 =>  inp_feat(487), I5 =>  inp_feat(336), I6 =>  inp_feat(370), I7 =>  inp_feat(496)); 
C_68_S_1_L_6_inst : LUT8 generic map(INIT => "1111101110100010111110111000000010101010100000101111111110001000001000001010000011000000100000000000000010000000100000000000000010011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_1_L_6_out, I0 =>  inp_feat(111), I1 =>  inp_feat(344), I2 =>  inp_feat(437), I3 =>  inp_feat(170), I4 =>  inp_feat(200), I5 =>  inp_feat(442), I6 =>  inp_feat(112), I7 =>  inp_feat(393)); 
C_68_S_1_L_7_inst : LUT8 generic map(INIT => "1010110011000000111111111111111101100100100000001110011011110010110001000000000011000100110000000000010001000000010001001100000010000000000000000000000000000000000000000000000000000000000000001000110000000000000001000000000000000100000000000000000000000000") port map( O =>C_68_S_1_L_7_out, I0 =>  inp_feat(297), I1 =>  inp_feat(234), I2 =>  inp_feat(49), I3 =>  inp_feat(370), I4 =>  inp_feat(265), I5 =>  inp_feat(372), I6 =>  inp_feat(145), I7 =>  inp_feat(393)); 
C_68_S_2_L_0_inst : LUT8 generic map(INIT => "1110110110101101000010001000110011001000100010001000000010001000100000010000000100000000000000000000000000000000000000000000000010001100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_2_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_68_S_2_L_1_inst : LUT8 generic map(INIT => "1110100010101010111000000000000010101000000000000000000000000000101010101010101000000000000000001010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001110100000001000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_2_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(372), I2 =>  inp_feat(442), I3 =>  inp_feat(347), I4 =>  inp_feat(393), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_68_S_2_L_2_inst : LUT8 generic map(INIT => "1010001000000000000000000000000010101010100000000010101000000000101000101100000010000000000000001000000010000000100000000000000011101010000000001000100000000000111011100000000000001010000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_68_S_2_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(278), I2 =>  inp_feat(442), I3 =>  inp_feat(393), I4 =>  inp_feat(241), I5 =>  inp_feat(283), I6 =>  inp_feat(89), I7 =>  inp_feat(336)); 
C_68_S_2_L_3_inst : LUT8 generic map(INIT => "1010000110101001100001011110011111111000101010100000000010100000111100011110000011000101110001011111001111100000000000001100001011110000101000000001010110100011111000001010000000000000101000001100000001000000000000010100000011110000110000000000000011000000") port map( O =>C_68_S_2_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(467), I2 =>  inp_feat(442), I3 =>  inp_feat(316), I4 =>  inp_feat(59), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(145)); 
C_68_S_2_L_4_inst : LUT8 generic map(INIT => "1110111000001100111011101000100011101100110001001100111000000000000010000000000000001000000000000000100000000000000010000000000010000000110000000000010000000000111111011100000010001110000000000000000000000000000000000000000000001000000000000000000000000000") port map( O =>C_68_S_2_L_4_out, I0 =>  inp_feat(372), I1 =>  inp_feat(442), I2 =>  inp_feat(180), I3 =>  inp_feat(312), I4 =>  inp_feat(65), I5 =>  inp_feat(478), I6 =>  inp_feat(44), I7 =>  inp_feat(195)); 
C_68_S_2_L_5_inst : LUT8 generic map(INIT => "0010111110101111101000101010001010100111101000001010000010000000101001101010001000000000000000001010001010100010000000000000000000101010001000000010001000000010101000000010000000000000000000001011110000100010000000000000000011100010001000100000000000000000") port map( O =>C_68_S_2_L_5_out, I0 =>  inp_feat(442), I1 =>  inp_feat(221), I2 =>  inp_feat(90), I3 =>  inp_feat(295), I4 =>  inp_feat(395), I5 =>  inp_feat(130), I6 =>  inp_feat(86), I7 =>  inp_feat(195)); 
C_68_S_2_L_6_inst : LUT8 generic map(INIT => "1110111111100000010000111100010011011101010011000100010111001100000000000000000000000000000000001000100000000000000000000000000000000000010001000000000011000100000000000000010000000000010001000000000000000000000000000100010000000000000001000000000001000100") port map( O =>C_68_S_2_L_6_out, I0 =>  inp_feat(351), I1 =>  inp_feat(106), I2 =>  inp_feat(440), I3 =>  inp_feat(471), I4 =>  inp_feat(111), I5 =>  inp_feat(462), I6 =>  inp_feat(168), I7 =>  inp_feat(393)); 
C_68_S_2_L_7_inst : LUT8 generic map(INIT => "1111111110110000000010100000000011110010000000001000101000000000111110101011000000000000000000000011000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000001010100000100000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_2_L_7_out, I0 =>  inp_feat(297), I1 =>  inp_feat(145), I2 =>  inp_feat(14), I3 =>  inp_feat(241), I4 =>  inp_feat(112), I5 =>  inp_feat(77), I6 =>  inp_feat(447), I7 =>  inp_feat(44)); 
C_68_S_3_L_0_inst : LUT8 generic map(INIT => "1110110110101101000010001000110011001000100010001000000010001000100000010000000100000000000000000000000000000000000000000000000010001100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_3_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_68_S_3_L_1_inst : LUT8 generic map(INIT => "1110100010101010111000000000000010101000000000000000000000000000101010101010101000000000000000001010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001110100000001000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_3_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(372), I2 =>  inp_feat(442), I3 =>  inp_feat(347), I4 =>  inp_feat(393), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_68_S_3_L_2_inst : LUT8 generic map(INIT => "1010001000000000000000000000000010101010100000000010101000000000101000101100000010000000000000001000000010000000100000000000000011101010000000001000100000000000111011100000000000001010000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_68_S_3_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(278), I2 =>  inp_feat(442), I3 =>  inp_feat(393), I4 =>  inp_feat(241), I5 =>  inp_feat(283), I6 =>  inp_feat(89), I7 =>  inp_feat(336)); 
C_68_S_3_L_3_inst : LUT8 generic map(INIT => "1011001110100000111001110010000111110010101100100010000000100000110001011100000011010101010001011111100111000000000000101100000011110000101000000011000100100011111000001010000000100000001000001100000001000000000000010100000011000000110000000100000011000000") port map( O =>C_68_S_3_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(9), I2 =>  inp_feat(442), I3 =>  inp_feat(111), I4 =>  inp_feat(59), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(145)); 
C_68_S_3_L_4_inst : LUT8 generic map(INIT => "0010111011001100110010001100010010001000100000000000000000000000101010101000100000001000100010001010000000000000001000000000000000101010111100001000100010100000101000000010000000000000000000001110101010001100000010000000110010101000000010000000100000000000") port map( O =>C_68_S_3_L_4_out, I0 =>  inp_feat(442), I1 =>  inp_feat(398), I2 =>  inp_feat(105), I3 =>  inp_feat(9), I4 =>  inp_feat(111), I5 =>  inp_feat(34), I6 =>  inp_feat(265), I7 =>  inp_feat(195)); 
C_68_S_3_L_5_inst : LUT8 generic map(INIT => "1111011011100110111111101110010000100000000000000010000001000000111111110010001011111111000000000000000000000000000000000000000000000000000000001111001000000000000000000000000000100000000000001111011100000000110111110000000000000000000000000000000000000000") port map( O =>C_68_S_3_L_5_out, I0 =>  inp_feat(336), I1 =>  inp_feat(221), I2 =>  inp_feat(312), I3 =>  inp_feat(209), I4 =>  inp_feat(478), I5 =>  inp_feat(44), I6 =>  inp_feat(171), I7 =>  inp_feat(195)); 
C_68_S_3_L_6_inst : LUT8 generic map(INIT => "1101011011110111011000101111001111000000011100110000000000000001101000001010000000000000000000000000000000000000000000000000000001000000000000000000000000000000110000001000000000000000000000001000000000000000000000000000000000000000001000000000000000000000") port map( O =>C_68_S_3_L_6_out, I0 =>  inp_feat(26), I1 =>  inp_feat(235), I2 =>  inp_feat(14), I3 =>  inp_feat(156), I4 =>  inp_feat(231), I5 =>  inp_feat(117), I6 =>  inp_feat(496), I7 =>  inp_feat(60)); 
C_68_S_3_L_7_inst : LUT8 generic map(INIT => "1111101111111110011111101111101100000000000000000001100000000000111111110001111110011100000111110000100000000000000110000000000001010010100100110011001100110011000000000000000000000000000000000011111100001011010100000000001100001000000000000000100000000000") port map( O =>C_68_S_3_L_7_out, I0 =>  inp_feat(480), I1 =>  inp_feat(108), I2 =>  inp_feat(336), I3 =>  inp_feat(180), I4 =>  inp_feat(437), I5 =>  inp_feat(168), I6 =>  inp_feat(462), I7 =>  inp_feat(158)); 
C_68_S_4_L_0_inst : LUT8 generic map(INIT => "1110110110101101000010001000110011001000100010001000000010001000100000010000000100000000000000000000000000000000000000000000000010001100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_4_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(44), I2 =>  inp_feat(82), I3 =>  inp_feat(363), I4 =>  inp_feat(442), I5 =>  inp_feat(347), I6 =>  inp_feat(393), I7 =>  inp_feat(117)); 
C_68_S_4_L_1_inst : LUT8 generic map(INIT => "1110100010101010111000000000000010101000000000000000000000000000101010101010101000000000000000001010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001110100000001000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_4_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(372), I2 =>  inp_feat(442), I3 =>  inp_feat(347), I4 =>  inp_feat(393), I5 =>  inp_feat(117), I6 =>  inp_feat(154), I7 =>  inp_feat(241)); 
C_68_S_4_L_2_inst : LUT8 generic map(INIT => "1010001000000000000000000000000010101010100000000010101000000000101000101100000010000000000000001000000010000000100000000000000011101010000000001000100000000000111011100000000000001010000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_68_S_4_L_2_out, I0 =>  inp_feat(168), I1 =>  inp_feat(278), I2 =>  inp_feat(442), I3 =>  inp_feat(393), I4 =>  inp_feat(241), I5 =>  inp_feat(283), I6 =>  inp_feat(89), I7 =>  inp_feat(336)); 
C_68_S_4_L_3_inst : LUT8 generic map(INIT => "1000001110100000111111011000000011101000101000101111100010000010111101000100000001110001111000001110000011000000111100111110000011000000111000101111000110100001000000001110000010000000100000000100000011000000000000010100000001000000110000000100000011000000") port map( O =>C_68_S_4_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(139), I2 =>  inp_feat(442), I3 =>  inp_feat(293), I4 =>  inp_feat(108), I5 =>  inp_feat(478), I6 =>  inp_feat(413), I7 =>  inp_feat(145)); 
C_68_S_4_L_4_inst : LUT8 generic map(INIT => "0100110011101101111110111110110011101000011011100010101000100000110000001110110100000000000011001000000011101100001000000000100010001000100010001000100010000000100010000000000000000000000000000000000010001000000000000000100010000000100010000000000000001000") port map( O =>C_68_S_4_L_4_out, I0 =>  inp_feat(33), I1 =>  inp_feat(442), I2 =>  inp_feat(172), I3 =>  inp_feat(478), I4 =>  inp_feat(329), I5 =>  inp_feat(390), I6 =>  inp_feat(424), I7 =>  inp_feat(34)); 
C_68_S_4_L_5_inst : LUT8 generic map(INIT => "1111111110101010101000001010100010100000100010000000000000000000011100100000000000100000001000100000000000000000000000000000000000100000001000000010000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000") port map( O =>C_68_S_4_L_5_out, I0 =>  inp_feat(499), I1 =>  inp_feat(452), I2 =>  inp_feat(434), I3 =>  inp_feat(145), I4 =>  inp_feat(14), I5 =>  inp_feat(241), I6 =>  inp_feat(112), I7 =>  inp_feat(44)); 
C_68_S_4_L_6_inst : LUT8 generic map(INIT => "1111110011111100011110001101010001010000010000000000000000000000110000000100000000000000000000000100000000000000000000000000000001010000100011000000100000001100010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_68_S_4_L_6_out, I0 =>  inp_feat(478), I1 =>  inp_feat(191), I2 =>  inp_feat(440), I3 =>  inp_feat(336), I4 =>  inp_feat(449), I5 =>  inp_feat(112), I6 =>  inp_feat(44), I7 =>  inp_feat(442)); 
C_68_S_4_L_7_inst : LUT8 generic map(INIT => "1111111100001111111101100000001011111111000001000011101000000000011111100000000011110010000000000010111000000000101010101000101011111100000000000100010000000000000001000000000000000100000000000011010000000000010101000000000000000100000000000000000000000000") port map( O =>C_68_S_4_L_7_out, I0 =>  inp_feat(331), I1 =>  inp_feat(494), I2 =>  inp_feat(180), I3 =>  inp_feat(349), I4 =>  inp_feat(7), I5 =>  inp_feat(364), I6 =>  inp_feat(372), I7 =>  inp_feat(49)); 
C_69_S_0_L_0_inst : LUT8 generic map(INIT => "1111111011101100111011111110000010001000100011001110111010001000010011101100110010001010101000000000100000001000000000000000000000000000000000000100100000000000100010001000100011001100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_0_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_69_S_0_L_1_inst : LUT8 generic map(INIT => "1111100011111101100000000010000010101000100000000000000000000000101010001111110100100000001000000000000000000000000000000000000000000000101010000000000000001000000000001000000000000000000000000000100010001000000000000000100000000000000000000000000000000000") port map( O =>C_69_S_0_L_1_out, I0 =>  inp_feat(389), I1 =>  inp_feat(347), I2 =>  inp_feat(102), I3 =>  inp_feat(336), I4 =>  inp_feat(349), I5 =>  inp_feat(276), I6 =>  inp_feat(295), I7 =>  inp_feat(370)); 
C_69_S_0_L_2_inst : LUT8 generic map(INIT => "0011001011111010101100101111001011101000110000001010000010001000110000001111000011110010111100101110100011000000010000000000000010001010110000001010000010100000101000001100000010000000000000000000000010000000000000000000000001000000110000000000000000000000") port map( O =>C_69_S_0_L_2_out, I0 =>  inp_feat(187), I1 =>  inp_feat(223), I2 =>  inp_feat(205), I3 =>  inp_feat(450), I4 =>  inp_feat(145), I5 =>  inp_feat(336), I6 =>  inp_feat(139), I7 =>  inp_feat(285)); 
C_69_S_0_L_3_inst : LUT8 generic map(INIT => "0111111110101011111011100111011110100000101000100000000000000111111110101011101101000000011100110000000010100010000000000000001111111100111100001111110001110000100000001010101010000000000000001100000000000000010000000000000010000000001000001000000010000000") port map( O =>C_69_S_0_L_3_out, I0 =>  inp_feat(285), I1 =>  inp_feat(26), I2 =>  inp_feat(450), I3 =>  inp_feat(54), I4 =>  inp_feat(452), I5 =>  inp_feat(279), I6 =>  inp_feat(388), I7 =>  inp_feat(301)); 
C_69_S_0_L_4_inst : LUT8 generic map(INIT => "1101101110000000000000001010101011111010000010001010001000001000001000000000000000000000000000000000100000000000000000000000000011111010100010001000000010001000111110100100000000100000000000001100100000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_0_L_4_out, I0 =>  inp_feat(277), I1 =>  inp_feat(183), I2 =>  inp_feat(413), I3 =>  inp_feat(488), I4 =>  inp_feat(442), I5 =>  inp_feat(86), I6 =>  inp_feat(503), I7 =>  inp_feat(82)); 
C_69_S_0_L_5_inst : LUT8 generic map(INIT => "1111110010111110000110101011101011111111100011101010101110101010111100001000110000001010000010101011101000001000101110101000101000000000000010000000000000000000000100001000100000000000000000101000000010000000000000000000000000110000100000000010000000000000") port map( O =>C_69_S_0_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(23), I2 =>  inp_feat(278), I3 =>  inp_feat(494), I4 =>  inp_feat(372), I5 =>  inp_feat(336), I6 =>  inp_feat(130), I7 =>  inp_feat(470)); 
C_69_S_0_L_6_inst : LUT8 generic map(INIT => "1111111000001100110111101110111000000000000000000100000000000000101010101010100011001100111010101000000000000000000000000000000010001010000010001000110000001000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_0_L_6_out, I0 =>  inp_feat(293), I1 =>  inp_feat(205), I2 =>  inp_feat(15), I3 =>  inp_feat(386), I4 =>  inp_feat(478), I5 =>  inp_feat(168), I6 =>  inp_feat(172), I7 =>  inp_feat(276)); 
C_69_S_0_L_7_inst : LUT8 generic map(INIT => "0111001010110000111111001111000000110000001100001111000010110000111110001011100010001000111100000010000000100000100000001111000011100000100000001111000011000000000000000000000010110000000000001100100000001000100000001000000000000000000000001000000010000000") port map( O =>C_69_S_0_L_7_out, I0 =>  inp_feat(69), I1 =>  inp_feat(46), I2 =>  inp_feat(442), I3 =>  inp_feat(321), I4 =>  inp_feat(478), I5 =>  inp_feat(411), I6 =>  inp_feat(171), I7 =>  inp_feat(295)); 
C_69_S_1_L_0_inst : LUT8 generic map(INIT => "1111111011101100111011111110000010001000100011001110111010001000010011101100110010001010101000000000100000001000000000000000000000000000000000000100100000000000100010001000100011001100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_1_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_69_S_1_L_1_inst : LUT8 generic map(INIT => "1111000011100100110000001100000011000000110011001100000011100000110001001100010011110000111100001010000001000100111100001111000000000000100000001000000010000000000000001000000000000000000000000000000000000000110010000000000000000000000000000000000000000000") port map( O =>C_69_S_1_L_1_out, I0 =>  inp_feat(280), I1 =>  inp_feat(150), I2 =>  inp_feat(44), I3 =>  inp_feat(450), I4 =>  inp_feat(249), I5 =>  inp_feat(244), I6 =>  inp_feat(277), I7 =>  inp_feat(370)); 
C_69_S_1_L_2_inst : LUT8 generic map(INIT => "0101110111111000110011001000100011001000000100001101111100000000010000001100000000000000000000000000110000000000000000000000000011111111110111000000000000000000110010101101000000000000000000001101110011001100000000000000000011001100010000000000110000000000") port map( O =>C_69_S_1_L_2_out, I0 =>  inp_feat(11), I1 =>  inp_feat(83), I2 =>  inp_feat(295), I3 =>  inp_feat(40), I4 =>  inp_feat(89), I5 =>  inp_feat(102), I6 =>  inp_feat(370), I7 =>  inp_feat(336)); 
C_69_S_1_L_3_inst : LUT8 generic map(INIT => "1111111000101010001010100010101000101110000000000000000000000000111110100000100010001010001010100000101000000000000000000000000011111010101010101011001000100000110010000000000000000000000000001111100000000000010100000000000011001000000000000000000000000000") port map( O =>C_69_S_1_L_3_out, I0 =>  inp_feat(442), I1 =>  inp_feat(478), I2 =>  inp_feat(26), I3 =>  inp_feat(117), I4 =>  inp_feat(23), I5 =>  inp_feat(241), I6 =>  inp_feat(388), I7 =>  inp_feat(302)); 
C_69_S_1_L_4_inst : LUT8 generic map(INIT => "0011101011110100111010001100111000100000000000001010100011101010000010000000000000100000000000000000000000000000000000000000000010100000100000001010000010000000101000001000000010100000000000000010000000000000111010000000000000000000000000001010101000000000") port map( O =>C_69_S_1_L_4_out, I0 =>  inp_feat(442), I1 =>  inp_feat(216), I2 =>  inp_feat(295), I3 =>  inp_feat(171), I4 =>  inp_feat(82), I5 =>  inp_feat(411), I6 =>  inp_feat(231), I7 =>  inp_feat(46)); 
C_69_S_1_L_5_inst : LUT8 generic map(INIT => "1000100011101011000000100000111010111111101111010000100010001100001010001000000000000000000000000010111000000000000000000000000011101010101010001000101010101110101000001011000000000000000000000000000010100000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_1_L_5_out, I0 =>  inp_feat(117), I1 =>  inp_feat(136), I2 =>  inp_feat(46), I3 =>  inp_feat(494), I4 =>  inp_feat(312), I5 =>  inp_feat(156), I6 =>  inp_feat(231), I7 =>  inp_feat(86)); 
C_69_S_1_L_6_inst : LUT8 generic map(INIT => "0010100000100000110110101000000011111101101000001000110000000000111110010000110111101100000011001010100110111000000011000000000010111011001000001010100010000000110111010000000000000000000000001011101000000000100000000000000000000000000000000000000000000000") port map( O =>C_69_S_1_L_6_out, I0 =>  inp_feat(370), I1 =>  inp_feat(43), I2 =>  inp_feat(483), I3 =>  inp_feat(470), I4 =>  inp_feat(82), I5 =>  inp_feat(145), I6 =>  inp_feat(302), I7 =>  inp_feat(7)); 
C_69_S_1_L_7_inst : LUT8 generic map(INIT => "0010110110100001000000011000101110011111100000000000000000000000111010001110111100000000010011111000101010000000000000000000000011111011111010011010101000101011111110110000000000101010000000001101000001101101000000000000001010001000000000000000000000000000") port map( O =>C_69_S_1_L_7_out, I0 =>  inp_feat(129), I1 =>  inp_feat(225), I2 =>  inp_feat(494), I3 =>  inp_feat(223), I4 =>  inp_feat(276), I5 =>  inp_feat(7), I6 =>  inp_feat(103), I7 =>  inp_feat(301)); 
C_69_S_2_L_0_inst : LUT8 generic map(INIT => "1111111011101100111011111110000010001000100011001110111010001000010011101100110010001010101000000000100000001000000000000000000000000000000000000100100000000000100010001000100011001100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_2_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_69_S_2_L_1_inst : LUT8 generic map(INIT => "0011001000010000111011111100001010100000000000001100000010000000101000001111000010111010111110001010000000000000000000000100000001111111011101010101011101011111101000100000000011000000100000000011000001110000000000000010000000100000000000000000000000000000") port map( O =>C_69_S_2_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(316), I2 =>  inp_feat(164), I3 =>  inp_feat(158), I4 =>  inp_feat(336), I5 =>  inp_feat(249), I6 =>  inp_feat(346), I7 =>  inp_feat(90)); 
C_69_S_2_L_2_inst : LUT8 generic map(INIT => "0010111011111011100011101000111111111100011100000000110000000000101011101011101100001111000011111111110011110000000001000000000011101100101000001110110010000000101010000000000000000000000000000000110000000000100010000000000000000000000000000000000000000000") port map( O =>C_69_S_2_L_2_out, I0 =>  inp_feat(215), I1 =>  inp_feat(89), I2 =>  inp_feat(82), I3 =>  inp_feat(450), I4 =>  inp_feat(283), I5 =>  inp_feat(359), I6 =>  inp_feat(149), I7 =>  inp_feat(302)); 
C_69_S_2_L_3_inst : LUT8 generic map(INIT => "1110101100101010111110101010101110001010000010001000000000000000110110100000000011110010101000001010000010100000101000001010000000111000000010000010001000000000101010111000001000000000000000001011101000100000101000101010000000100000101000001010000000100000") port map( O =>C_69_S_2_L_3_out, I0 =>  inp_feat(117), I1 =>  inp_feat(108), I2 =>  inp_feat(180), I3 =>  inp_feat(468), I4 =>  inp_feat(228), I5 =>  inp_feat(462), I6 =>  inp_feat(121), I7 =>  inp_feat(297)); 
C_69_S_2_L_4_inst : LUT8 generic map(INIT => "0010101110101111101010000000111011111111110011110110111011101110111111011000111110100000100000001111000000000000000000000000000000000000000000010000000000000000100010000000000000000000000000001000111100001111000000000000000010000000000000000000000000000000") port map( O =>C_69_S_2_L_4_out, I0 =>  inp_feat(269), I1 =>  inp_feat(149), I2 =>  inp_feat(336), I3 =>  inp_feat(130), I4 =>  inp_feat(256), I5 =>  inp_feat(478), I6 =>  inp_feat(305), I7 =>  inp_feat(258)); 
C_69_S_2_L_5_inst : LUT8 generic map(INIT => "0110110110110000111101111111101011011110110011101111111110001111111101001011000011010000111100001100000010000000010000000000000000000000000000001100000000000000000000000000000000000000000000001100010000000000110000000000000000000000000000000000000000000000") port map( O =>C_69_S_2_L_5_out, I0 =>  inp_feat(331), I1 =>  inp_feat(33), I2 =>  inp_feat(378), I3 =>  inp_feat(145), I4 =>  inp_feat(478), I5 =>  inp_feat(329), I6 =>  inp_feat(388), I7 =>  inp_feat(258)); 
C_69_S_2_L_6_inst : LUT8 generic map(INIT => "1110111111110111111011111000000010000000101100011100110010000000111101111111110111111010000000000000000000000001000000000000000011000000100000001100000000000000000000001000000000001100100000000100000000000000110000000000000000000000000000000000000000000000") port map( O =>C_69_S_2_L_6_out, I0 =>  inp_feat(359), I1 =>  inp_feat(153), I2 =>  inp_feat(183), I3 =>  inp_feat(61), I4 =>  inp_feat(149), I5 =>  inp_feat(326), I6 =>  inp_feat(499), I7 =>  inp_feat(503)); 
C_69_S_2_L_7_inst : LUT8 generic map(INIT => "0110111111111100001000000010100011100100111011001110000011100000101111110000010010101010000000001111010100000000000000000000000001100100101000000000000000100000111000001010000010100000101000001111111100000000101010000000000011110101000000000000000000000000") port map( O =>C_69_S_2_L_7_out, I0 =>  inp_feat(154), I1 =>  inp_feat(457), I2 =>  inp_feat(388), I3 =>  inp_feat(336), I4 =>  inp_feat(83), I5 =>  inp_feat(329), I6 =>  inp_feat(89), I7 =>  inp_feat(37)); 
C_69_S_3_L_0_inst : LUT8 generic map(INIT => "1111111011101100111011111110000010001000100011001110111010001000010011101100110010001010101000000000100000001000000000000000000000000000000000000100100000000000100010001000100011001100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_3_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_69_S_3_L_1_inst : LUT8 generic map(INIT => "0011001000010000111011111100001010100000000000001100000010000000101000001111000010111010111110001010000000000000000000000100000001111111011101010101011101011111101000100000000011000000100000000011000001110000000000000010000000100000000000000000000000000000") port map( O =>C_69_S_3_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(316), I2 =>  inp_feat(164), I3 =>  inp_feat(158), I4 =>  inp_feat(336), I5 =>  inp_feat(249), I6 =>  inp_feat(346), I7 =>  inp_feat(90)); 
C_69_S_3_L_2_inst : LUT8 generic map(INIT => "0010101010110011100010101010001010111011111100110000101100000010111110001011000000001000000000001000000010110000000000000000000010111011111100001000100010000000100110101011000010001000000000001010100000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_3_L_2_out, I0 =>  inp_feat(117), I1 =>  inp_feat(484), I2 =>  inp_feat(82), I3 =>  inp_feat(450), I4 =>  inp_feat(283), I5 =>  inp_feat(145), I6 =>  inp_feat(359), I7 =>  inp_feat(302)); 
C_69_S_3_L_3_inst : LUT8 generic map(INIT => "1111111000100010111111100011000001001100000000001111100000110000101010100000000010001000000000001000100000000000100010001000000000100110000001000000000000000000000000000000000001000000000000001010011100000000101000000000000010000000000000001000100010000000") port map( O =>C_69_S_3_L_3_out, I0 =>  inp_feat(145), I1 =>  inp_feat(82), I2 =>  inp_feat(436), I3 =>  inp_feat(503), I4 =>  inp_feat(46), I5 =>  inp_feat(37), I6 =>  inp_feat(86), I7 =>  inp_feat(370)); 
C_69_S_3_L_4_inst : LUT8 generic map(INIT => "1101100111100001110000001000000001000000000010000000000000000000110111111101110110000000100000001100100110101110100000000000100001000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000000011000000000010000000000000000000") port map( O =>C_69_S_3_L_4_out, I0 =>  inp_feat(46), I1 =>  inp_feat(132), I2 =>  inp_feat(408), I3 =>  inp_feat(336), I4 =>  inp_feat(442), I5 =>  inp_feat(474), I6 =>  inp_feat(478), I7 =>  inp_feat(117)); 
C_69_S_3_L_5_inst : LUT8 generic map(INIT => "0111111111101010101100001110000011010000100000000010000010100000111010100110101010100000110000001100000010000000100000001100000001100010010000000000100000000000000000000000000000000000000000001110111011000000100010001100000000000000010000001000000001000000") port map( O =>C_69_S_3_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(89), I2 =>  inp_feat(230), I3 =>  inp_feat(265), I4 =>  inp_feat(333), I5 =>  inp_feat(321), I6 =>  inp_feat(171), I7 =>  inp_feat(347)); 
C_69_S_3_L_6_inst : LUT8 generic map(INIT => "1111011111011011111100111111101110101111101000100010000010100000110000101011000001011011101110001000001010010010000000000000000001110001000000000000000010000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_3_L_6_out, I0 =>  inp_feat(295), I1 =>  inp_feat(478), I2 =>  inp_feat(427), I3 =>  inp_feat(301), I4 =>  inp_feat(380), I5 =>  inp_feat(117), I6 =>  inp_feat(113), I7 =>  inp_feat(168)); 
C_69_S_3_L_7_inst : LUT8 generic map(INIT => "0010000011000000110000001100000010101110101011001000000000000000111110001100000010000000100000000010000000000000100000000000000011110010010000001100000001000000101110100000000010000000000000001111000000000000101000000000000000100000000000000000000000000000") port map( O =>C_69_S_3_L_7_out, I0 =>  inp_feat(83), I1 =>  inp_feat(307), I2 =>  inp_feat(442), I3 =>  inp_feat(405), I4 =>  inp_feat(223), I5 =>  inp_feat(302), I6 =>  inp_feat(291), I7 =>  inp_feat(7)); 
C_69_S_4_L_0_inst : LUT8 generic map(INIT => "1111111011101100111011111110000010001000100011001110111010001000010011101100110010001010101000000000100000001000000000000000000000000000000000000100100000000000100010001000100011001100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_4_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_69_S_4_L_1_inst : LUT8 generic map(INIT => "0011001000010000111011111100001010100000000000001100000010000000101000001111000010111010111110001010000000000000000000000100000001111111011101010101011101011111101000100000000011000000100000000011000001110000000000000010000000100000000000000000000000000000") port map( O =>C_69_S_4_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(316), I2 =>  inp_feat(164), I3 =>  inp_feat(158), I4 =>  inp_feat(336), I5 =>  inp_feat(249), I6 =>  inp_feat(346), I7 =>  inp_feat(90)); 
C_69_S_4_L_2_inst : LUT8 generic map(INIT => "0010101010110011100010101010001010111011111100110000101100000010111110001011000000001000000000001000000010110000000000000000000010111011111100001000100010000000100110101011000010001000000000001010100000000000000000000000000000000000000000000000000000000000") port map( O =>C_69_S_4_L_2_out, I0 =>  inp_feat(117), I1 =>  inp_feat(484), I2 =>  inp_feat(82), I3 =>  inp_feat(450), I4 =>  inp_feat(283), I5 =>  inp_feat(145), I6 =>  inp_feat(359), I7 =>  inp_feat(302)); 
C_69_S_4_L_3_inst : LUT8 generic map(INIT => "1111111000100010111111100011000001001100000000001111100000110000101010100000000010001000000000001000100000000000100010001000000000100110000001000000000000000000000000000000000001000000000000001010011100000000101000000000000010000000000000001000100010000000") port map( O =>C_69_S_4_L_3_out, I0 =>  inp_feat(145), I1 =>  inp_feat(82), I2 =>  inp_feat(436), I3 =>  inp_feat(503), I4 =>  inp_feat(46), I5 =>  inp_feat(37), I6 =>  inp_feat(86), I7 =>  inp_feat(370)); 
C_69_S_4_L_4_inst : LUT8 generic map(INIT => "1101110010111100110001001100110001000000110011000000000000000000111111111011111110000000000010001101001011011101100000000001001001001100000000000000000000000000000000000000000000000000000000001111100000000000000000000000000001000000010100000000000000000000") port map( O =>C_69_S_4_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(411), I2 =>  inp_feat(413), I3 =>  inp_feat(336), I4 =>  inp_feat(442), I5 =>  inp_feat(474), I6 =>  inp_feat(478), I7 =>  inp_feat(117)); 
C_69_S_4_L_5_inst : LUT8 generic map(INIT => "1101110011011010010011001000100011111100101011001000100010001100110101001101000011001100000000001100000010001000000000001000100000001000100010101000000000000000000000000000000000000000000000001000000000000000100000000000000010000000000000001000000000000000") port map( O =>C_69_S_4_L_5_out, I0 =>  inp_feat(121), I1 =>  inp_feat(132), I2 =>  inp_feat(149), I3 =>  inp_feat(336), I4 =>  inp_feat(183), I5 =>  inp_feat(249), I6 =>  inp_feat(285), I7 =>  inp_feat(164)); 
C_69_S_4_L_6_inst : LUT8 generic map(INIT => "0111111011111000111110101010100000100000100000000010000000000000111011100100000000101010000000000010000000000000001000100000000000001100110000000000000000000000000000000000000000000000000000001100110011000000000000000000000010001000000000000000000000000000") port map( O =>C_69_S_4_L_6_out, I0 =>  inp_feat(508), I1 =>  inp_feat(26), I2 =>  inp_feat(228), I3 =>  inp_feat(64), I4 =>  inp_feat(121), I5 =>  inp_feat(349), I6 =>  inp_feat(485), I7 =>  inp_feat(347)); 
C_69_S_4_L_7_inst : LUT8 generic map(INIT => "1111001011110010101110111010101000100010101000001010101110101010111110001100000011011110100010100000001010000000000010101000101010010000000000001000100000000000101000100000000010101010000000000011000000000000000000100000000000000000000000000000001000000000") port map( O =>C_69_S_4_L_7_out, I0 =>  inp_feat(442), I1 =>  inp_feat(336), I2 =>  inp_feat(195), I3 =>  inp_feat(179), I4 =>  inp_feat(478), I5 =>  inp_feat(107), I6 =>  inp_feat(78), I7 =>  inp_feat(83)); 
C_70_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(86), I2 =>  inp_feat(187), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_70_S_0_L_1_inst : LUT8 generic map(INIT => "1100100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_1_out, I0 =>  inp_feat(511), I1 =>  inp_feat(200), I2 =>  inp_feat(276), I3 =>  inp_feat(7), I4 =>  inp_feat(450), I5 =>  inp_feat(249), I6 =>  inp_feat(330), I7 =>  inp_feat(329)); 
C_70_S_0_L_2_inst : LUT8 generic map(INIT => "0010000000000000000000000000000010100000101000000000000000000000000010000000001000000000000100000000000000000000000000000000000010100000100010000100000000000000101000001010000001010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_2_out, I0 =>  inp_feat(234), I1 =>  inp_feat(347), I2 =>  inp_feat(352), I3 =>  inp_feat(437), I4 =>  inp_feat(15), I5 =>  inp_feat(205), I6 =>  inp_feat(336), I7 =>  inp_feat(370)); 
C_70_S_0_L_3_inst : LUT8 generic map(INIT => "1101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_3_out, I0 =>  inp_feat(499), I1 =>  inp_feat(38), I2 =>  inp_feat(238), I3 =>  inp_feat(491), I4 =>  inp_feat(86), I5 =>  inp_feat(26), I6 =>  inp_feat(82), I7 =>  inp_feat(388)); 
C_70_S_0_L_4_inst : LUT8 generic map(INIT => "1000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000") port map( O =>C_70_S_0_L_4_out, I0 =>  inp_feat(7), I1 =>  inp_feat(316), I2 =>  inp_feat(26), I3 =>  inp_feat(82), I4 =>  inp_feat(121), I5 =>  inp_feat(283), I6 =>  inp_feat(210), I7 =>  inp_feat(414)); 
C_70_S_0_L_5_inst : LUT8 generic map(INIT => "0001000000000000000000000000000011001000000000000000000001000000100000000000000000000000100000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_5_out, I0 =>  inp_feat(136), I1 =>  inp_feat(218), I2 =>  inp_feat(220), I3 =>  inp_feat(511), I4 =>  inp_feat(478), I5 =>  inp_feat(398), I6 =>  inp_feat(499), I7 =>  inp_feat(81)); 
C_70_S_0_L_6_inst : LUT8 generic map(INIT => "1000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_6_out, I0 =>  inp_feat(139), I1 =>  inp_feat(484), I2 =>  inp_feat(1), I3 =>  inp_feat(149), I4 =>  inp_feat(424), I5 =>  inp_feat(403), I6 =>  inp_feat(151), I7 =>  inp_feat(347)); 
C_70_S_0_L_7_inst : LUT8 generic map(INIT => "1101000011000000000000001100000010000000110000000000000000000000001000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_0_L_7_out, I0 =>  inp_feat(493), I1 =>  inp_feat(71), I2 =>  inp_feat(457), I3 =>  inp_feat(132), I4 =>  inp_feat(336), I5 =>  inp_feat(268), I6 =>  inp_feat(34), I7 =>  inp_feat(8)); 
C_70_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_1_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(86), I2 =>  inp_feat(187), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_70_S_1_L_1_inst : LUT8 generic map(INIT => "1101110000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_1_L_1_out, I0 =>  inp_feat(499), I1 =>  inp_feat(336), I2 =>  inp_feat(276), I3 =>  inp_feat(7), I4 =>  inp_feat(450), I5 =>  inp_feat(249), I6 =>  inp_feat(330), I7 =>  inp_feat(329)); 
C_70_S_1_L_2_inst : LUT8 generic map(INIT => "0000001000000000000000000100000001100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000110000000000000000000000100000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_1_L_2_out, I0 =>  inp_feat(347), I1 =>  inp_feat(210), I2 =>  inp_feat(283), I3 =>  inp_feat(107), I4 =>  inp_feat(108), I5 =>  inp_feat(294), I6 =>  inp_feat(316), I7 =>  inp_feat(398)); 
C_70_S_1_L_3_inst : LUT8 generic map(INIT => "1010000010100010000000000000000000000000100000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_1_L_3_out, I0 =>  inp_feat(53), I1 =>  inp_feat(158), I2 =>  inp_feat(64), I3 =>  inp_feat(100), I4 =>  inp_feat(291), I5 =>  inp_feat(302), I6 =>  inp_feat(462), I7 =>  inp_feat(149)); 
C_70_S_1_L_4_inst : LUT8 generic map(INIT => "1100000110000000000000001000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000010000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_1_L_4_out, I0 =>  inp_feat(136), I1 =>  inp_feat(504), I2 =>  inp_feat(413), I3 =>  inp_feat(354), I4 =>  inp_feat(302), I5 =>  inp_feat(82), I6 =>  inp_feat(347), I7 =>  inp_feat(164)); 
C_70_S_1_L_5_inst : LUT8 generic map(INIT => "1000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000") port map( O =>C_70_S_1_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(413), I2 =>  inp_feat(475), I3 =>  inp_feat(145), I4 =>  inp_feat(238), I5 =>  inp_feat(462), I6 =>  inp_feat(352), I7 =>  inp_feat(49)); 
C_70_S_1_L_6_inst : LUT8 generic map(INIT => "0010001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000010010000000000001000100010000000000000000000000000000000000000000000000000000000100000000000000000001000") port map( O =>C_70_S_1_L_6_out, I0 =>  inp_feat(173), I1 =>  inp_feat(443), I2 =>  inp_feat(148), I3 =>  inp_feat(190), I4 =>  inp_feat(336), I5 =>  inp_feat(234), I6 =>  inp_feat(478), I7 =>  inp_feat(499)); 
C_70_S_1_L_7_inst : LUT8 generic map(INIT => "0010000010101010101000001010000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_1_L_7_out, I0 =>  inp_feat(82), I1 =>  inp_feat(338), I2 =>  inp_feat(336), I3 =>  inp_feat(347), I4 =>  inp_feat(201), I5 =>  inp_feat(131), I6 =>  inp_feat(283), I7 =>  inp_feat(388)); 
C_70_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_2_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(86), I2 =>  inp_feat(187), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_70_S_2_L_1_inst : LUT8 generic map(INIT => "1101110000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_2_L_1_out, I0 =>  inp_feat(499), I1 =>  inp_feat(336), I2 =>  inp_feat(276), I3 =>  inp_feat(7), I4 =>  inp_feat(450), I5 =>  inp_feat(249), I6 =>  inp_feat(330), I7 =>  inp_feat(329)); 
C_70_S_2_L_2_inst : LUT8 generic map(INIT => "0000001010000000000000000000100010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_2_L_2_out, I0 =>  inp_feat(330), I1 =>  inp_feat(412), I2 =>  inp_feat(357), I3 =>  inp_feat(148), I4 =>  inp_feat(108), I5 =>  inp_feat(294), I6 =>  inp_feat(316), I7 =>  inp_feat(398)); 
C_70_S_2_L_3_inst : LUT8 generic map(INIT => "1110000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_2_L_3_out, I0 =>  inp_feat(131), I1 =>  inp_feat(357), I2 =>  inp_feat(491), I3 =>  inp_feat(82), I4 =>  inp_feat(40), I5 =>  inp_feat(387), I6 =>  inp_feat(462), I7 =>  inp_feat(149)); 
C_70_S_2_L_4_inst : LUT8 generic map(INIT => "1000000000000000000000000000000011000000000000001100000000000000101000000000000010000000000000001100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100000") port map( O =>C_70_S_2_L_4_out, I0 =>  inp_feat(98), I1 =>  inp_feat(357), I2 =>  inp_feat(151), I3 =>  inp_feat(388), I4 =>  inp_feat(396), I5 =>  inp_feat(132), I6 =>  inp_feat(338), I7 =>  inp_feat(336)); 
C_70_S_2_L_5_inst : LUT8 generic map(INIT => "1000000000100000100000000000000000000000000000000000000010000000000000001000000010100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000") port map( O =>C_70_S_2_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(53), I2 =>  inp_feat(180), I3 =>  inp_feat(34), I4 =>  inp_feat(386), I5 =>  inp_feat(478), I6 =>  inp_feat(107), I7 =>  inp_feat(256)); 
C_70_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000010000000000000010000000010000000000000000000000100000000000000000000000000000001100000000000000000000000000000000010000000000000000000000000000101100000000000000000000000000000000000100000000000000000000000010100000000000000000000000000000") port map( O =>C_70_S_2_L_6_out, I0 =>  inp_feat(183), I1 =>  inp_feat(406), I2 =>  inp_feat(64), I3 =>  inp_feat(109), I4 =>  inp_feat(90), I5 =>  inp_feat(442), I6 =>  inp_feat(148), I7 =>  inp_feat(110)); 
C_70_S_2_L_7_inst : LUT8 generic map(INIT => "1000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_2_L_7_out, I0 =>  inp_feat(86), I1 =>  inp_feat(146), I2 =>  inp_feat(145), I3 =>  inp_feat(204), I4 =>  inp_feat(302), I5 =>  inp_feat(291), I6 =>  inp_feat(215), I7 =>  inp_feat(13)); 
C_70_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(86), I2 =>  inp_feat(187), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_70_S_3_L_1_inst : LUT8 generic map(INIT => "1001100100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_1_out, I0 =>  inp_feat(150), I1 =>  inp_feat(462), I2 =>  inp_feat(11), I3 =>  inp_feat(200), I4 =>  inp_feat(450), I5 =>  inp_feat(249), I6 =>  inp_feat(330), I7 =>  inp_feat(329)); 
C_70_S_3_L_2_inst : LUT8 generic map(INIT => "0000000000001001100010000000100000000000100000000000000010001000000001000000110000000000000000001000000000100000000000000000000000000000000000000000100010001000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_2_out, I0 =>  inp_feat(171), I1 =>  inp_feat(331), I2 =>  inp_feat(212), I3 =>  inp_feat(158), I4 =>  inp_feat(125), I5 =>  inp_feat(326), I6 =>  inp_feat(111), I7 =>  inp_feat(98)); 
C_70_S_3_L_3_inst : LUT8 generic map(INIT => "0101000010000000110100000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_3_out, I0 =>  inp_feat(44), I1 =>  inp_feat(58), I2 =>  inp_feat(283), I3 =>  inp_feat(371), I4 =>  inp_feat(437), I5 =>  inp_feat(352), I6 =>  inp_feat(149), I7 =>  inp_feat(98)); 
C_70_S_3_L_4_inst : LUT8 generic map(INIT => "1000100000000000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_4_out, I0 =>  inp_feat(215), I1 =>  inp_feat(363), I2 =>  inp_feat(148), I3 =>  inp_feat(145), I4 =>  inp_feat(117), I5 =>  inp_feat(316), I6 =>  inp_feat(453), I7 =>  inp_feat(130)); 
C_70_S_3_L_5_inst : LUT8 generic map(INIT => "1000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_5_out, I0 =>  inp_feat(185), I1 =>  inp_feat(17), I2 =>  inp_feat(478), I3 =>  inp_feat(19), I4 =>  inp_feat(283), I5 =>  inp_feat(295), I6 =>  inp_feat(131), I7 =>  inp_feat(84)); 
C_70_S_3_L_6_inst : LUT8 generic map(INIT => "0000100000100000100000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000001000000100000000110010000000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_6_out, I0 =>  inp_feat(352), I1 =>  inp_feat(372), I2 =>  inp_feat(136), I3 =>  inp_feat(265), I4 =>  inp_feat(499), I5 =>  inp_feat(413), I6 =>  inp_feat(462), I7 =>  inp_feat(474)); 
C_70_S_3_L_7_inst : LUT8 generic map(INIT => "0100001011000000000000001000000011011000000010000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_3_L_7_out, I0 =>  inp_feat(347), I1 =>  inp_feat(336), I2 =>  inp_feat(197), I3 =>  inp_feat(111), I4 =>  inp_feat(93), I5 =>  inp_feat(409), I6 =>  inp_feat(125), I7 =>  inp_feat(220)); 
C_70_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_0_out, I0 =>  inp_feat(336), I1 =>  inp_feat(86), I2 =>  inp_feat(187), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_70_S_4_L_1_inst : LUT8 generic map(INIT => "1001100100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_1_out, I0 =>  inp_feat(150), I1 =>  inp_feat(462), I2 =>  inp_feat(11), I3 =>  inp_feat(200), I4 =>  inp_feat(450), I5 =>  inp_feat(249), I6 =>  inp_feat(330), I7 =>  inp_feat(329)); 
C_70_S_4_L_2_inst : LUT8 generic map(INIT => "1000000000000000010100010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000010000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_2_out, I0 =>  inp_feat(49), I1 =>  inp_feat(405), I2 =>  inp_feat(357), I3 =>  inp_feat(316), I4 =>  inp_feat(158), I5 =>  inp_feat(221), I6 =>  inp_feat(265), I7 =>  inp_feat(98)); 
C_70_S_4_L_3_inst : LUT8 generic map(INIT => "1010001000100010000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_3_out, I0 =>  inp_feat(450), I1 =>  inp_feat(158), I2 =>  inp_feat(331), I3 =>  inp_feat(265), I4 =>  inp_feat(302), I5 =>  inp_feat(120), I6 =>  inp_feat(90), I7 =>  inp_feat(82)); 
C_70_S_4_L_4_inst : LUT8 generic map(INIT => "0000000011100000000000000000000000010000000000000000000000000000111100100111001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_4_out, I0 =>  inp_feat(347), I1 =>  inp_feat(107), I2 =>  inp_feat(249), I3 =>  inp_feat(205), I4 =>  inp_feat(475), I5 =>  inp_feat(336), I6 =>  inp_feat(370), I7 =>  inp_feat(352)); 
C_70_S_4_L_5_inst : LUT8 generic map(INIT => "1000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010001000000000000000000000000000100010001000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(272), I2 =>  inp_feat(94), I3 =>  inp_feat(420), I4 =>  inp_feat(145), I5 =>  inp_feat(303), I6 =>  inp_feat(352), I7 =>  inp_feat(470)); 
C_70_S_4_L_6_inst : LUT8 generic map(INIT => "0001000000000000111100000000000000000000000000001000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000001101000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_6_out, I0 =>  inp_feat(186), I1 =>  inp_feat(505), I2 =>  inp_feat(456), I3 =>  inp_feat(149), I4 =>  inp_feat(326), I5 =>  inp_feat(352), I6 =>  inp_feat(425), I7 =>  inp_feat(164)); 
C_70_S_4_L_7_inst : LUT8 generic map(INIT => "0000100000000000100000000000000011000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_70_S_4_L_7_out, I0 =>  inp_feat(82), I1 =>  inp_feat(286), I2 =>  inp_feat(111), I3 =>  inp_feat(108), I4 =>  inp_feat(425), I5 =>  inp_feat(164), I6 =>  inp_feat(302), I7 =>  inp_feat(380)); 
C_71_S_0_L_0_inst : LUT8 generic map(INIT => "1111111011011000111010101010000010001100100010001010101010001000010011101000110010001010101000000000110000001000000000000000000000000000000000001000100000000000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_0_L_0_out, I0 =>  inp_feat(459), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_71_S_0_L_1_inst : LUT8 generic map(INIT => "1110101011110111111000001000000000111111110100001110110010000000100010001101000010000000000000001001110011010100110011001000000000110010011100110000000000000000000100000101000000001100000000000011000001010000000000000000000011111001010100000000100000000000") port map( O =>C_71_S_0_L_1_out, I0 =>  inp_feat(362), I1 =>  inp_feat(0), I2 =>  inp_feat(318), I3 =>  inp_feat(462), I4 =>  inp_feat(279), I5 =>  inp_feat(437), I6 =>  inp_feat(295), I7 =>  inp_feat(370)); 
C_71_S_0_L_2_inst : LUT8 generic map(INIT => "0110001010010000001100100011001110111011000010100101101100001011111100001111000011100000000000001100000010000000110000000000000011110000000000001111000111111111111111100000001000111111101010111100000000000000111000000000000000000000000000000000000000000000") port map( O =>C_71_S_0_L_2_out, I0 =>  inp_feat(469), I1 =>  inp_feat(336), I2 =>  inp_feat(193), I3 =>  inp_feat(187), I4 =>  inp_feat(437), I5 =>  inp_feat(331), I6 =>  inp_feat(450), I7 =>  inp_feat(154)); 
C_71_S_0_L_3_inst : LUT8 generic map(INIT => "0011110011111001111010101110000011001100110111011000000011010001111000001110100010100000101000000100010000000000000000000000000001000000110001000000000000000000110000000000000110000000000000001110000010001000100000000000000011000000000000001100000000000000") port map( O =>C_71_S_0_L_3_out, I0 =>  inp_feat(336), I1 =>  inp_feat(129), I2 =>  inp_feat(25), I3 =>  inp_feat(478), I4 =>  inp_feat(145), I5 =>  inp_feat(82), I6 =>  inp_feat(286), I7 =>  inp_feat(442)); 
C_71_S_0_L_4_inst : LUT8 generic map(INIT => "0111111111111110011101101100000000110110110001001110011011010100111111001000100000000000000000001100000000000000110000000100000000010100000000000000000000000000000000000000000000000000010000001111100010001000010000001100000000000000000000001100000001000000") port map( O =>C_71_S_0_L_4_out, I0 =>  inp_feat(478), I1 =>  inp_feat(223), I2 =>  inp_feat(228), I3 =>  inp_feat(336), I4 =>  inp_feat(387), I5 =>  inp_feat(297), I6 =>  inp_feat(30), I7 =>  inp_feat(148)); 
C_71_S_0_L_5_inst : LUT8 generic map(INIT => "1010111110111010111011110000001000001101111111111100111100001111111110001111100010101100000000000101000011110000110010000000000000000000000000001100000000000000000000000000000001000100000000001000000000000000000000000000000000000000000100000000000000000000") port map( O =>C_71_S_0_L_5_out, I0 =>  inp_feat(493), I1 =>  inp_feat(11), I2 =>  inp_feat(249), I3 =>  inp_feat(86), I4 =>  inp_feat(178), I5 =>  inp_feat(107), I6 =>  inp_feat(78), I7 =>  inp_feat(503)); 
C_71_S_0_L_6_inst : LUT8 generic map(INIT => "0010110000111111001000110010111100111100001111110010001000111011111110000000000011110010000100000000100100000000001100100000000011111111011101111010000000100001101010000010000000100000001000001010101000000010000000000000000000001000000000000000000000000000") port map( O =>C_71_S_0_L_6_out, I0 =>  inp_feat(107), I1 =>  inp_feat(478), I2 =>  inp_feat(329), I3 =>  inp_feat(143), I4 =>  inp_feat(167), I5 =>  inp_feat(111), I6 =>  inp_feat(220), I7 =>  inp_feat(420)); 
C_71_S_0_L_7_inst : LUT8 generic map(INIT => "0111001111110110011100101010111000101010111011100010001010101110111000101111111011111000111011100010000011101110000000001000111011110011111000010000000000000000100000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_0_L_7_out, I0 =>  inp_feat(302), I1 =>  inp_feat(145), I2 =>  inp_feat(107), I3 =>  inp_feat(478), I4 =>  inp_feat(468), I5 =>  inp_feat(493), I6 =>  inp_feat(413), I7 =>  inp_feat(17)); 
C_71_S_1_L_0_inst : LUT8 generic map(INIT => "1111111011011000111010101010000010001100100010001010101010001000010011101000110010001010101000000000110000001000000000000000000000000000000000001000100000000000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_1_L_0_out, I0 =>  inp_feat(459), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_71_S_1_L_1_inst : LUT8 generic map(INIT => "1100101010001111111011111010111111101111101011110000000010101111000000110000001100000000001100111100111110101011000000000000111100001010000000011100111100000011100011111000111110000100000011111000000000000000000000000000000010001000100010100000000000000000") port map( O =>C_71_S_1_L_1_out, I0 =>  inp_feat(411), I1 =>  inp_feat(195), I2 =>  inp_feat(478), I3 =>  inp_feat(462), I4 =>  inp_feat(378), I5 =>  inp_feat(108), I6 =>  inp_feat(94), I7 =>  inp_feat(111)); 
C_71_S_1_L_2_inst : LUT8 generic map(INIT => "0101110110001010111111110000101011111111000010001111101100000000010011110000101001001111000011001110111100001010000011110000000011000000000010001110101000001010010100000000000001010000000000000100000001001100000000000000000000000000000000000000000000000000") port map( O =>C_71_S_1_L_2_out, I0 =>  inp_feat(154), I1 =>  inp_feat(380), I2 =>  inp_feat(478), I3 =>  inp_feat(136), I4 =>  inp_feat(109), I5 =>  inp_feat(413), I6 =>  inp_feat(86), I7 =>  inp_feat(456)); 
C_71_S_1_L_3_inst : LUT8 generic map(INIT => "0010000011110000111000001110010011100100101000000010000000000000111111011111010101000100010101001110000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000001000100000000000000010000000000010001000000000000000000000000000") port map( O =>C_71_S_1_L_3_out, I0 =>  inp_feat(336), I1 =>  inp_feat(17), I2 =>  inp_feat(503), I3 =>  inp_feat(420), I4 =>  inp_feat(322), I5 =>  inp_feat(145), I6 =>  inp_feat(82), I7 =>  inp_feat(231)); 
C_71_S_1_L_4_inst : LUT8 generic map(INIT => "0110101011001000110010001000100011111000110010001000100010000000111111101010000010111111101010001110101000000000100011000000000000000000000000000000000010001000000000000000000000000000000000000000001000000000000000001000100000000010000000000000000000000000") port map( O =>C_71_S_1_L_4_out, I0 =>  inp_feat(357), I1 =>  inp_feat(62), I2 =>  inp_feat(249), I3 =>  inp_feat(316), I4 =>  inp_feat(221), I5 =>  inp_feat(388), I6 =>  inp_feat(180), I7 =>  inp_feat(231)); 
C_71_S_1_L_5_inst : LUT8 generic map(INIT => "0111001010100010111110001110100001000000000000000100010000000000111100001010000001010000101010100000000000000000000000000000000000100010101010101010111011101110000000000010101000000000000000000001000010000000101111001000111000000000000000000000000000000000") port map( O =>C_71_S_1_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(86), I2 =>  inp_feat(166), I3 =>  inp_feat(494), I4 =>  inp_feat(329), I5 =>  inp_feat(231), I6 =>  inp_feat(153), I7 =>  inp_feat(11)); 
C_71_S_1_L_6_inst : LUT8 generic map(INIT => "1011111111001001000000000101000011001111110101010000000111010001101001001000000010000000000000001100010010000000101110011000000000001100100000000000000000000000110011011000100010000000000000001100110010000000101000000000000011001100100000001010000000000000") port map( O =>C_71_S_1_L_6_out, I0 =>  inp_feat(427), I1 =>  inp_feat(347), I2 =>  inp_feat(7), I3 =>  inp_feat(103), I4 =>  inp_feat(458), I5 =>  inp_feat(494), I6 =>  inp_feat(329), I7 =>  inp_feat(11)); 
C_71_S_1_L_7_inst : LUT8 generic map(INIT => "1111111010001000011110101011101011001000100001000000000000000000110011000010101000001000101010101000110000000000000000000000000010001000000010000000100000000000000010001000100000000000000000001000100000001010000010000000111000001000000000000000000000000000") port map( O =>C_71_S_1_L_7_out, I0 =>  inp_feat(442), I1 =>  inp_feat(148), I2 =>  inp_feat(478), I3 =>  inp_feat(49), I4 =>  inp_feat(111), I5 =>  inp_feat(43), I6 =>  inp_feat(424), I7 =>  inp_feat(100)); 
C_71_S_2_L_0_inst : LUT8 generic map(INIT => "1111111011011000111010101010000010001100100010001010101010001000010011101000110010001010101000000000110000001000000000000000000000000000000000001000100000000000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_2_L_0_out, I0 =>  inp_feat(459), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_71_S_2_L_1_inst : LUT8 generic map(INIT => "0000111011101000111111111010001011001011110010100000000010000000100010001100100011111111111000000000000011000000000000001100000011101000110000001010100000000000110010000100000000000000000000001000100010001000100000000000000000000000000000000000000000000000") port map( O =>C_71_S_2_L_1_out, I0 =>  inp_feat(470), I1 =>  inp_feat(499), I2 =>  inp_feat(7), I3 =>  inp_feat(154), I4 =>  inp_feat(82), I5 =>  inp_feat(227), I6 =>  inp_feat(295), I7 =>  inp_feat(291)); 
C_71_S_2_L_2_inst : LUT8 generic map(INIT => "1110111101110110111000100010001001000111010011101000101110001011111010000000010000000000000000001100000000000100100000000000000001010011011100000000000000100000110000110000100010000000000000001111101101010000000000000000000011000000000000000000000000000000") port map( O =>C_71_S_2_L_2_out, I0 =>  inp_feat(90), I1 =>  inp_feat(462), I2 =>  inp_feat(62), I3 =>  inp_feat(158), I4 =>  inp_feat(322), I5 =>  inp_feat(327), I6 =>  inp_feat(145), I7 =>  inp_feat(293)); 
C_71_S_2_L_3_inst : LUT8 generic map(INIT => "0111010011100110000000001100010011100000110000001111000001000000111010001100110000000000110011001110000001000100101000000100000011101100100011001100000011001100101000000000000010100000000000001100010010001100110000001100110010100000000000001010000000000000") port map( O =>C_71_S_2_L_3_out, I0 =>  inp_feat(333), I1 =>  inp_feat(305), I2 =>  inp_feat(158), I3 =>  inp_feat(336), I4 =>  inp_feat(505), I5 =>  inp_feat(103), I6 =>  inp_feat(302), I7 =>  inp_feat(450)); 
C_71_S_2_L_4_inst : LUT8 generic map(INIT => "0010111011111001101010111111011110110000111100001000000011010100000000001000000010000000100000000000000010000000000000001000000011101000100000011100101011111111111100001111000011000000110001000000000000000000100000001000000000000000000000001100000010000000") port map( O =>C_71_S_2_L_4_out, I0 =>  inp_feat(256), I1 =>  inp_feat(130), I2 =>  inp_feat(287), I3 =>  inp_feat(478), I4 =>  inp_feat(82), I5 =>  inp_feat(99), I6 =>  inp_feat(231), I7 =>  inp_feat(329)); 
C_71_S_2_L_5_inst : LUT8 generic map(INIT => "0111110111011101111000000110110011111001001000001010100000100000000010000000100000000000000000001111000000000000001000000000000000000000010000001100000001110000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000") port map( O =>C_71_S_2_L_5_out, I0 =>  inp_feat(46), I1 =>  inp_feat(180), I2 =>  inp_feat(260), I3 =>  inp_feat(357), I4 =>  inp_feat(336), I5 =>  inp_feat(9), I6 =>  inp_feat(148), I7 =>  inp_feat(101)); 
C_71_S_2_L_6_inst : LUT8 generic map(INIT => "1111101000000000110110101000001011011100110000001101100011001000011110101101000011111010111100100000000001000000010100000100000000001000000000001101100001000000100000001000000011010000110000000000000000000000000000000000000000000000000000000101000000000000") port map( O =>C_71_S_2_L_6_out, I0 =>  inp_feat(180), I1 =>  inp_feat(295), I2 =>  inp_feat(127), I3 =>  inp_feat(347), I4 =>  inp_feat(336), I5 =>  inp_feat(64), I6 =>  inp_feat(437), I7 =>  inp_feat(101)); 
C_71_S_2_L_7_inst : LUT8 generic map(INIT => "1111110111010100110000001000000011110111000001001111001111000000010111010010000011011010101010000000111100100000000001011010101011001101010101011000000010000000001011111010111000001011101010100000100111101100000001001010101000000111101010100000011110101010") port map( O =>C_71_S_2_L_7_out, I0 =>  inp_feat(478), I1 =>  inp_feat(107), I2 =>  inp_feat(0), I3 =>  inp_feat(54), I4 =>  inp_feat(228), I5 =>  inp_feat(99), I6 =>  inp_feat(303), I7 =>  inp_feat(323)); 
C_71_S_3_L_0_inst : LUT8 generic map(INIT => "1111111011011000111010101010000010001100100010001010101010001000010011101000110010001010101000000000110000001000000000000000000000000000000000001000100000000000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_3_L_0_out, I0 =>  inp_feat(459), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_71_S_3_L_1_inst : LUT8 generic map(INIT => "0111000011101000111000101110000011110000111100000000000010100000100000001010100011100000111000000000000010100000000000001010000011110010110000001111001000000000010000001000000000000000000000001110000010000000010000100000000000000000000000000000000000000000") port map( O =>C_71_S_3_L_1_out, I0 =>  inp_feat(48), I1 =>  inp_feat(316), I2 =>  inp_feat(231), I3 =>  inp_feat(154), I4 =>  inp_feat(82), I5 =>  inp_feat(227), I6 =>  inp_feat(295), I7 =>  inp_feat(291)); 
C_71_S_3_L_2_inst : LUT8 generic map(INIT => "1111011101111111001100001101000011010001000100001101010111010001111001000000000011100000000000001000000000000000101000000000000001110000010100000000000000000000011100000111000000000000000000001100000000000000110011000000000010000000000000000000000000000000") port map( O =>C_71_S_3_L_2_out, I0 =>  inp_feat(478), I1 =>  inp_feat(329), I2 =>  inp_feat(148), I3 =>  inp_feat(304), I4 =>  inp_feat(68), I5 =>  inp_feat(322), I6 =>  inp_feat(209), I7 =>  inp_feat(232)); 
C_71_S_3_L_3_inst : LUT8 generic map(INIT => "1101111101100010011110100010101001110101011000000110010100000000000010100000000000101010000000100001000100000000001000010000000011001110110011101100111011001110101011000100110000000000010000000000100000001100000011100000111000001000000001000000000000000000") port map( O =>C_71_S_3_L_3_out, I0 =>  inp_feat(81), I1 =>  inp_feat(472), I2 =>  inp_feat(248), I3 =>  inp_feat(411), I4 =>  inp_feat(280), I5 =>  inp_feat(11), I6 =>  inp_feat(111), I7 =>  inp_feat(249)); 
C_71_S_3_L_4_inst : LUT8 generic map(INIT => "1100111100010101101011100000000011001101000000000000100000000000111011101110010010101111101000001110111010000000000010110010000011001100010001000000000000000000010010000100000000000000000000001100110011001100000000000000000011001100100011000000000000000000") port map( O =>C_71_S_3_L_4_out, I0 =>  inp_feat(23), I1 =>  inp_feat(111), I2 =>  inp_feat(265), I3 =>  inp_feat(83), I4 =>  inp_feat(327), I5 =>  inp_feat(222), I6 =>  inp_feat(81), I7 =>  inp_feat(400)); 
C_71_S_3_L_5_inst : LUT8 generic map(INIT => "1100100010000100110110001100100001000100110010000000000000000000010100000000000011111100100000000100000000000000000000001000000011011110010011000000111110001010010011101100110000001010100010001111111000000000010011101000100000000010000000000000100010000000") port map( O =>C_71_S_3_L_5_out, I0 =>  inp_feat(121), I1 =>  inp_feat(470), I2 =>  inp_feat(483), I3 =>  inp_feat(80), I4 =>  inp_feat(336), I5 =>  inp_feat(111), I6 =>  inp_feat(212), I7 =>  inp_feat(108)); 
C_71_S_3_L_6_inst : LUT8 generic map(INIT => "1011011011101010111110101110100101001001000110111111111111011111111100000111000011110000011100000010000000000000011000000010000001000000110000000000000011100000000000000000000000000000000000000100000000000000010000000010000000000000000000000000000000000000") port map( O =>C_71_S_3_L_6_out, I0 =>  inp_feat(472), I1 =>  inp_feat(265), I2 =>  inp_feat(312), I3 =>  inp_feat(221), I4 =>  inp_feat(478), I5 =>  inp_feat(386), I6 =>  inp_feat(155), I7 =>  inp_feat(148)); 
C_71_S_3_L_7_inst : LUT8 generic map(INIT => "0101110101011111110101010101010110000101000000001001100100000000110100001101000011010000100100001000000000000000100000001000000011101101000011001010110100000101110011110000000000001111000010011000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_71_S_3_L_7_out, I0 =>  inp_feat(329), I1 =>  inp_feat(187), I2 =>  inp_feat(46), I3 =>  inp_feat(41), I4 =>  inp_feat(149), I5 =>  inp_feat(501), I6 =>  inp_feat(220), I7 =>  inp_feat(305)); 
C_71_S_4_L_0_inst : LUT8 generic map(INIT => "1111111011011000111010101010000010001100100010001010101010001000010011101000110010001010101000000000110000001000000000000000000000000000000000001000100000000000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_4_L_0_out, I0 =>  inp_feat(459), I1 =>  inp_feat(83), I2 =>  inp_feat(478), I3 =>  inp_feat(82), I4 =>  inp_feat(260), I5 =>  inp_feat(484), I6 =>  inp_feat(499), I7 =>  inp_feat(117)); 
C_71_S_4_L_1_inst : LUT8 generic map(INIT => "0111111000001000111011100010000011111111000000000000101000000000100010100000100011101110000000000000101000000000000010100000000011111100001000001111000000100000010010000000000000000000000000001110100000000000010000000010000000000000000000000000000000000000") port map( O =>C_71_S_4_L_1_out, I0 =>  inp_feat(48), I1 =>  inp_feat(316), I2 =>  inp_feat(154), I3 =>  inp_feat(231), I4 =>  inp_feat(82), I5 =>  inp_feat(227), I6 =>  inp_feat(295), I7 =>  inp_feat(291)); 
C_71_S_4_L_2_inst : LUT8 generic map(INIT => "1111001011100000110100001100000011111111111111111110000101010000100000000100000001000000110000000000000011001100010000001100010011110110111100000100000011001000010101101111111100000010010001010000000000000000010000000100000001000000000000000100000001000000") port map( O =>C_71_S_4_L_2_out, I0 =>  inp_feat(413), I1 =>  inp_feat(273), I2 =>  inp_feat(499), I3 =>  inp_feat(265), I4 =>  inp_feat(437), I5 =>  inp_feat(331), I6 =>  inp_feat(68), I7 =>  inp_feat(232)); 
C_71_S_4_L_3_inst : LUT8 generic map(INIT => "1011101111101010101010101010100000000000101000000010000010101000000000001000000010101010100000000000000001000000000000001000100011101010110010100000100000001000100000001000100000001000000010001000100000000000101011101000110000000000000000000000100000001000") port map( O =>C_71_S_4_L_3_out, I0 =>  inp_feat(117), I1 =>  inp_feat(439), I2 =>  inp_feat(167), I3 =>  inp_feat(467), I4 =>  inp_feat(336), I5 =>  inp_feat(186), I6 =>  inp_feat(370), I7 =>  inp_feat(249)); 
C_71_S_4_L_4_inst : LUT8 generic map(INIT => "1101111101000011111111001100000011111111000000001111111110000000110011010000110011010000110000001101110100001100101100111000000000001000000000001010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_71_S_4_L_4_out, I0 =>  inp_feat(467), I1 =>  inp_feat(386), I2 =>  inp_feat(81), I3 =>  inp_feat(111), I4 =>  inp_feat(457), I5 =>  inp_feat(303), I6 =>  inp_feat(483), I7 =>  inp_feat(258)); 
C_71_S_4_L_5_inst : LUT8 generic map(INIT => "1101111011001101111111001000110000001000100000001101100000000000110010101000000011001000000011001100100000000000110010000000000010001000100010001011101000001100000000000000000000000000000000001010101000000000101011100000110000000000000000000000000000000000") port map( O =>C_71_S_4_L_5_out, I0 =>  inp_feat(411), I1 =>  inp_feat(470), I2 =>  inp_feat(336), I3 =>  inp_feat(333), I4 =>  inp_feat(180), I5 =>  inp_feat(326), I6 =>  inp_feat(200), I7 =>  inp_feat(440)); 
C_71_S_4_L_6_inst : LUT8 generic map(INIT => "0101110111111000110000001111010111101010000010000111101100110110110000001111010000000000001100000000000000000000000000000000010011001010101011101000000000000010110010000000000010001010000000001010000011101110100010001010111000000000000000000000000000000000") port map( O =>C_71_S_4_L_6_out, I0 =>  inp_feat(7), I1 =>  inp_feat(297), I2 =>  inp_feat(505), I3 =>  inp_feat(333), I4 =>  inp_feat(321), I5 =>  inp_feat(46), I6 =>  inp_feat(153), I7 =>  inp_feat(82)); 
C_71_S_4_L_7_inst : LUT8 generic map(INIT => "1011111010001110111111101011101000111110000000101111111000111010111011001010101001101100001010101000101000000000000000000000000000000000000000000000100000000000000010000000000000000000000000001000100010001010001010000010101000001000000000000000000000000000") port map( O =>C_71_S_4_L_7_out, I0 =>  inp_feat(347), I1 =>  inp_feat(265), I2 =>  inp_feat(494), I3 =>  inp_feat(411), I4 =>  inp_feat(302), I5 =>  inp_feat(437), I6 =>  inp_feat(484), I7 =>  inp_feat(117)); 
C_72_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000010000000000000000000000000000000000000000001000000000100000000000000010000010000000000000000000000000000000000000000000000000000100000110000100000001000000010001001010000010000000100000000000000010000000100000000000000000000000") port map( O =>C_72_S_0_L_0_out, I0 =>  inp_feat(217), I1 =>  inp_feat(210), I2 =>  inp_feat(98), I3 =>  inp_feat(502), I4 =>  inp_feat(429), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_72_S_0_L_1_inst : LUT8 generic map(INIT => "1010000000100000010000000000000011110101000000000010000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_0_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(331), I2 =>  inp_feat(98), I3 =>  inp_feat(494), I4 =>  inp_feat(366), I5 =>  inp_feat(502), I6 =>  inp_feat(492), I7 =>  inp_feat(388)); 
C_72_S_0_L_2_inst : LUT8 generic map(INIT => "0010000110101110111100001111000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_0_L_2_out, I0 =>  inp_feat(365), I1 =>  inp_feat(155), I2 =>  inp_feat(375), I3 =>  inp_feat(6), I4 =>  inp_feat(265), I5 =>  inp_feat(422), I6 =>  inp_feat(219), I7 =>  inp_feat(420)); 
C_72_S_0_L_3_inst : LUT8 generic map(INIT => "0011000010110000110000000101000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000001000001110100001100000001010000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_0_L_3_out, I0 =>  inp_feat(80), I1 =>  inp_feat(451), I2 =>  inp_feat(58), I3 =>  inp_feat(381), I4 =>  inp_feat(505), I5 =>  inp_feat(349), I6 =>  inp_feat(227), I7 =>  inp_feat(65)); 
C_72_S_0_L_4_inst : LUT8 generic map(INIT => "1101000011010110000000000000000001100000010110000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_0_L_4_out, I0 =>  inp_feat(220), I1 =>  inp_feat(161), I2 =>  inp_feat(494), I3 =>  inp_feat(82), I4 =>  inp_feat(415), I5 =>  inp_feat(65), I6 =>  inp_feat(328), I7 =>  inp_feat(350)); 
C_72_S_0_L_5_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000001000101000000000000000000000000000001000000000000010000000000000101010100000000010000010000010100000000000000000000000000000000000001010000000011010000000001000001010000000000000100000000000000000101000010000") port map( O =>C_72_S_0_L_5_out, I0 =>  inp_feat(420), I1 =>  inp_feat(238), I2 =>  inp_feat(167), I3 =>  inp_feat(102), I4 =>  inp_feat(281), I5 =>  inp_feat(323), I6 =>  inp_feat(437), I7 =>  inp_feat(413)); 
C_72_S_0_L_6_inst : LUT8 generic map(INIT => "0010010010000000101010100010001000000010000000001010000100000000000000000000000010100000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_0_L_6_out, I0 =>  inp_feat(494), I1 =>  inp_feat(357), I2 =>  inp_feat(437), I3 =>  inp_feat(102), I4 =>  inp_feat(281), I5 =>  inp_feat(85), I6 =>  inp_feat(137), I7 =>  inp_feat(276)); 
C_72_S_0_L_7_inst : LUT8 generic map(INIT => "1101011000000000111100010000001000000000000000001010000000000000100001000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000010000000000000000000000") port map( O =>C_72_S_0_L_7_out, I0 =>  inp_feat(206), I1 =>  inp_feat(469), I2 =>  inp_feat(388), I3 =>  inp_feat(504), I4 =>  inp_feat(281), I5 =>  inp_feat(91), I6 =>  inp_feat(21), I7 =>  inp_feat(494)); 
C_72_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000010000000000000000000000000000000000000000001000000000100000000000000010000010000000000000000000000000000000000000000000000000000100000110000100000001000000010001001010000010000000100000000000000010000000100000000000000000000000") port map( O =>C_72_S_1_L_0_out, I0 =>  inp_feat(217), I1 =>  inp_feat(210), I2 =>  inp_feat(98), I3 =>  inp_feat(502), I4 =>  inp_feat(429), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_72_S_1_L_1_inst : LUT8 generic map(INIT => "1010000000100000010000000000000011110101000000000010000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_1_L_1_out, I0 =>  inp_feat(100), I1 =>  inp_feat(331), I2 =>  inp_feat(98), I3 =>  inp_feat(494), I4 =>  inp_feat(366), I5 =>  inp_feat(502), I6 =>  inp_feat(492), I7 =>  inp_feat(388)); 
C_72_S_1_L_2_inst : LUT8 generic map(INIT => "1010001010001000101000000100100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_1_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(280), I2 =>  inp_feat(58), I3 =>  inp_feat(375), I4 =>  inp_feat(65), I5 =>  inp_feat(422), I6 =>  inp_feat(219), I7 =>  inp_feat(420)); 
C_72_S_1_L_3_inst : LUT8 generic map(INIT => "0000110001000100000000001101010000000100010000000000000011000101000000000000010000000000100000001000000000000000110000001100010001000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010100000000000000010000000000000") port map( O =>C_72_S_1_L_3_out, I0 =>  inp_feat(281), I1 =>  inp_feat(494), I2 =>  inp_feat(155), I3 =>  inp_feat(323), I4 =>  inp_feat(238), I5 =>  inp_feat(413), I6 =>  inp_feat(74), I7 =>  inp_feat(500)); 
C_72_S_1_L_4_inst : LUT8 generic map(INIT => "0000000000011100000000000000000000011100001010100100000001101000000000000000000000000000000000000000010000000000000000000000000000001010100010100000000000000000000010000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_1_L_4_out, I0 =>  inp_feat(509), I1 =>  inp_feat(182), I2 =>  inp_feat(265), I3 =>  inp_feat(6), I4 =>  inp_feat(388), I5 =>  inp_feat(65), I6 =>  inp_feat(276), I7 =>  inp_feat(268)); 
C_72_S_1_L_5_inst : LUT8 generic map(INIT => "0100110000000010001011000000000000000000010000000000000000000000000000000000000000000000000001010000000000000000000000000000000000101110101000001000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_1_L_5_out, I0 =>  inp_feat(65), I1 =>  inp_feat(115), I2 =>  inp_feat(80), I3 =>  inp_feat(241), I4 =>  inp_feat(282), I5 =>  inp_feat(349), I6 =>  inp_feat(504), I7 =>  inp_feat(167)); 
C_72_S_1_L_6_inst : LUT8 generic map(INIT => "0001000100010010001010100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011110100000000011011001100000000000000000000000000000000000000001001000000000000100100000000000010000000000000000000000000000000") port map( O =>C_72_S_1_L_6_out, I0 =>  inp_feat(105), I1 =>  inp_feat(237), I2 =>  inp_feat(352), I3 =>  inp_feat(123), I4 =>  inp_feat(505), I5 =>  inp_feat(400), I6 =>  inp_feat(85), I7 =>  inp_feat(381)); 
C_72_S_1_L_7_inst : LUT8 generic map(INIT => "1100101011000000000000001100000000000000000000000000000011000000000000000100000001000000000000000000000000000000000000000000000000001001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_1_L_7_out, I0 =>  inp_feat(352), I1 =>  inp_feat(494), I2 =>  inp_feat(286), I3 =>  inp_feat(47), I4 =>  inp_feat(3), I5 =>  inp_feat(422), I6 =>  inp_feat(396), I7 =>  inp_feat(240)); 
C_72_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000010000000000000000000000000000000000000000001000000000100000000000000010000010000000000000000000000000000000000000000000000000000100000110000100000001000000010001001010000010000000100000000000000010000000100000000000000000000000") port map( O =>C_72_S_2_L_0_out, I0 =>  inp_feat(217), I1 =>  inp_feat(210), I2 =>  inp_feat(98), I3 =>  inp_feat(502), I4 =>  inp_feat(429), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_72_S_2_L_1_inst : LUT8 generic map(INIT => "1101110000000000100000000000000011011100000000000100000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_2_L_1_out, I0 =>  inp_feat(87), I1 =>  inp_feat(429), I2 =>  inp_feat(11), I3 =>  inp_feat(330), I4 =>  inp_feat(366), I5 =>  inp_feat(502), I6 =>  inp_feat(492), I7 =>  inp_feat(388)); 
C_72_S_2_L_2_inst : LUT8 generic map(INIT => "1000110011001000000000001000000001001000110011000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_2_L_2_out, I0 =>  inp_feat(353), I1 =>  inp_feat(504), I2 =>  inp_feat(19), I3 =>  inp_feat(80), I4 =>  inp_feat(316), I5 =>  inp_feat(193), I6 =>  inp_feat(399), I7 =>  inp_feat(494)); 
C_72_S_2_L_3_inst : LUT8 generic map(INIT => "0000100000000000000000000000100000001000100010001000110000001000000000000000000000000000000000000000000000000000000000000000000000001010100010000000000000000000000010001000101010110000000000000000000000000000000000000000000000000000100000000000000000000000") port map( O =>C_72_S_2_L_3_out, I0 =>  inp_feat(477), I1 =>  inp_feat(494), I2 =>  inp_feat(469), I3 =>  inp_feat(406), I4 =>  inp_feat(476), I5 =>  inp_feat(206), I6 =>  inp_feat(345), I7 =>  inp_feat(65)); 
C_72_S_2_L_4_inst : LUT8 generic map(INIT => "0000000110010110000000000000000011100100111101000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_2_L_4_out, I0 =>  inp_feat(65), I1 =>  inp_feat(182), I2 =>  inp_feat(509), I3 =>  inp_feat(6), I4 =>  inp_feat(422), I5 =>  inp_feat(265), I6 =>  inp_feat(316), I7 =>  inp_feat(219)); 
C_72_S_2_L_5_inst : LUT8 generic map(INIT => "0000010100110000111000000000000100000000000000001111001100000000000000000000000000000001000000000000000000000000111000000000000010110000100000000000000000000000010000000000000011100000000000000000000000000000000000000000000011000000000000000100000000000000") port map( O =>C_72_S_2_L_5_out, I0 =>  inp_feat(297), I1 =>  inp_feat(65), I2 =>  inp_feat(280), I3 =>  inp_feat(494), I4 =>  inp_feat(455), I5 =>  inp_feat(167), I6 =>  inp_feat(350), I7 =>  inp_feat(74)); 
C_72_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000000000100010000000100010010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000001100100000000000100000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_2_L_6_out, I0 =>  inp_feat(280), I1 =>  inp_feat(232), I2 =>  inp_feat(368), I3 =>  inp_feat(58), I4 =>  inp_feat(172), I5 =>  inp_feat(241), I6 =>  inp_feat(276), I7 =>  inp_feat(502)); 
C_72_S_2_L_7_inst : LUT8 generic map(INIT => "1000001010000010000000000011010000000000001000000000000000000000000000110010001000001000110000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000001011001000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_2_L_7_out, I0 =>  inp_feat(178), I1 =>  inp_feat(357), I2 =>  inp_feat(116), I3 =>  inp_feat(331), I4 =>  inp_feat(375), I5 =>  inp_feat(422), I6 =>  inp_feat(467), I7 =>  inp_feat(350)); 
C_72_S_3_L_0_inst : LUT8 generic map(INIT => "0000000010000000000000000000000100000000000000000000000000000000000010001000100011000100010011000000000000000000000000000000000000000010110010110000100000001001000000000000000000000000100000000000000000000000110011011000111100001000000000000000000000000000") port map( O =>C_72_S_3_L_0_out, I0 =>  inp_feat(109), I1 =>  inp_feat(193), I2 =>  inp_feat(6), I3 =>  inp_feat(469), I4 =>  inp_feat(406), I5 =>  inp_feat(494), I6 =>  inp_feat(438), I7 =>  inp_feat(206)); 
C_72_S_3_L_1_inst : LUT8 generic map(INIT => "1010100000000000000000000000000000000000000000000000000000000000101000000010000000000000000000000110000000000000000100000000000010101000000100000010000000100000000000000000000000000000000000001010000000010000000000000000000001000000000000000001000001000000") port map( O =>C_72_S_3_L_1_out, I0 =>  inp_feat(494), I1 =>  inp_feat(238), I2 =>  inp_feat(345), I3 =>  inp_feat(420), I4 =>  inp_feat(178), I5 =>  inp_feat(363), I6 =>  inp_feat(382), I7 =>  inp_feat(65)); 
C_72_S_3_L_2_inst : LUT8 generic map(INIT => "0010000000000000000000000000000000000010100000000000000000000000000000100000000000000000000000000000001000000000000000000000000010100000000000000000000000000000101010100000000000000000000000000000000000001000100000000000000000000000000000000000000000000000") port map( O =>C_72_S_3_L_2_out, I0 =>  inp_feat(309), I1 =>  inp_feat(505), I2 =>  inp_feat(280), I3 =>  inp_feat(58), I4 =>  inp_feat(471), I5 =>  inp_feat(409), I6 =>  inp_feat(349), I7 =>  inp_feat(502)); 
C_72_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000110100000001000100000000000000000000000000010001010011110000100110000000000110011100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000") port map( O =>C_72_S_3_L_3_out, I0 =>  inp_feat(468), I1 =>  inp_feat(280), I2 =>  inp_feat(65), I3 =>  inp_feat(180), I4 =>  inp_feat(324), I5 =>  inp_feat(350), I6 =>  inp_feat(6), I7 =>  inp_feat(328)); 
C_72_S_3_L_4_inst : LUT8 generic map(INIT => "0100100000001010010010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011000000111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_3_L_4_out, I0 =>  inp_feat(348), I1 =>  inp_feat(494), I2 =>  inp_feat(375), I3 =>  inp_feat(31), I4 =>  inp_feat(247), I5 =>  inp_feat(422), I6 =>  inp_feat(276), I7 =>  inp_feat(293)); 
C_72_S_3_L_5_inst : LUT8 generic map(INIT => "0010000000100000000000001000000011000000101000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011100001110000001100000000000000000000000000000101000000000000000100000000000000000000000000000") port map( O =>C_72_S_3_L_5_out, I0 =>  inp_feat(509), I1 =>  inp_feat(74), I2 =>  inp_feat(52), I3 =>  inp_feat(256), I4 =>  inp_feat(494), I5 =>  inp_feat(339), I6 =>  inp_feat(498), I7 =>  inp_feat(380)); 
C_72_S_3_L_6_inst : LUT8 generic map(INIT => "0011100110000000101100000000000000000000000000000000000000100000000100000000000011010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000") port map( O =>C_72_S_3_L_6_out, I0 =>  inp_feat(80), I1 =>  inp_feat(65), I2 =>  inp_feat(375), I3 =>  inp_feat(345), I4 =>  inp_feat(338), I5 =>  inp_feat(422), I6 =>  inp_feat(167), I7 =>  inp_feat(396)); 
C_72_S_3_L_7_inst : LUT8 generic map(INIT => "0000000100010101000000000001000010100000001100000000000000000000000000000100000000000000000000000000000000000000000000000000000001010001010100000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_3_L_7_out, I0 =>  inp_feat(80), I1 =>  inp_feat(206), I2 =>  inp_feat(41), I3 =>  inp_feat(65), I4 =>  inp_feat(477), I5 =>  inp_feat(83), I6 =>  inp_feat(366), I7 =>  inp_feat(101)); 
C_72_S_4_L_0_inst : LUT8 generic map(INIT => "0000000010000000000000000000000100000000000000000000000000000000000010001000100011000100010011000000000000000000000000000000000000000010110010110000100000001001000000000000000000000000100000000000000000000000110011011000111100001000000000000000000000000000") port map( O =>C_72_S_4_L_0_out, I0 =>  inp_feat(109), I1 =>  inp_feat(193), I2 =>  inp_feat(6), I3 =>  inp_feat(469), I4 =>  inp_feat(406), I5 =>  inp_feat(494), I6 =>  inp_feat(438), I7 =>  inp_feat(206)); 
C_72_S_4_L_1_inst : LUT8 generic map(INIT => "1110001000010000000000000000000000000000000000000000000000000000101000010011000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_4_L_1_out, I0 =>  inp_feat(286), I1 =>  inp_feat(238), I2 =>  inp_feat(60), I3 =>  inp_feat(178), I4 =>  inp_feat(219), I5 =>  inp_feat(227), I6 =>  inp_feat(65), I7 =>  inp_feat(349)); 
C_72_S_4_L_2_inst : LUT8 generic map(INIT => "0110000000000000000000000000000000000000000000000000000000000000010000000000000011000000010000000100000001000000001000000000000011000000000000000000000000000000000000000000000000000000000000001110000010000010010000000000000000000000000000100000000000000000") port map( O =>C_72_S_4_L_2_out, I0 =>  inp_feat(256), I1 =>  inp_feat(30), I2 =>  inp_feat(504), I3 =>  inp_feat(494), I4 =>  inp_feat(280), I5 =>  inp_feat(420), I6 =>  inp_feat(65), I7 =>  inp_feat(380)); 
C_72_S_4_L_3_inst : LUT8 generic map(INIT => "1100101000000000010010000000000010101010001000000000101000000000000000000000000010000000000000001010101000000000000010000000001000000000000000000000000000000000000001000000000000000000000000000000000000000100100000000000000000001000001000000000000000000000") port map( O =>C_72_S_4_L_3_out, I0 =>  inp_feat(232), I1 =>  inp_feat(329), I2 =>  inp_feat(256), I3 =>  inp_feat(494), I4 =>  inp_feat(280), I5 =>  inp_feat(206), I6 =>  inp_feat(21), I7 =>  inp_feat(420)); 
C_72_S_4_L_4_inst : LUT8 generic map(INIT => "0100010001000100010001000100010000000100010101001101110001000100000001000000000000000000000000010000101000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000") port map( O =>C_72_S_4_L_4_out, I0 =>  inp_feat(80), I1 =>  inp_feat(494), I2 =>  inp_feat(105), I3 =>  inp_feat(65), I4 =>  inp_feat(62), I5 =>  inp_feat(390), I6 =>  inp_feat(247), I7 =>  inp_feat(422)); 
C_72_S_4_L_5_inst : LUT8 generic map(INIT => "0110000010000000000000001000100000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000010000000101000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_4_L_5_out, I0 =>  inp_feat(53), I1 =>  inp_feat(355), I2 =>  inp_feat(491), I3 =>  inp_feat(319), I4 =>  inp_feat(397), I5 =>  inp_feat(422), I6 =>  inp_feat(276), I7 =>  inp_feat(268)); 
C_72_S_4_L_6_inst : LUT8 generic map(INIT => "0111000100000000000000000000000000100000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000011010000000000000010001000100000000000000000000010000000000000001000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_72_S_4_L_6_out, I0 =>  inp_feat(206), I1 =>  inp_feat(129), I2 =>  inp_feat(494), I3 =>  inp_feat(504), I4 =>  inp_feat(366), I5 =>  inp_feat(349), I6 =>  inp_feat(405), I7 =>  inp_feat(427)); 
C_72_S_4_L_7_inst : LUT8 generic map(INIT => "0000011000000000000000010000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010000000000000000010000010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_72_S_4_L_7_out, I0 =>  inp_feat(316), I1 =>  inp_feat(429), I2 =>  inp_feat(80), I3 =>  inp_feat(88), I4 =>  inp_feat(102), I5 =>  inp_feat(459), I6 =>  inp_feat(422), I7 =>  inp_feat(167)); 
C_73_S_0_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000001000001000000000000000000000000000000000001000000000000000000000000010100000000000001010000000000000101000000000000000100000000000001010000000000000") port map( O =>C_73_S_0_L_0_out, I0 =>  inp_feat(128), I1 =>  inp_feat(351), I2 =>  inp_feat(178), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_73_S_0_L_1_inst : LUT8 generic map(INIT => "0000000100000000000010000000000000000100000000000100010000000000000000000000000000000000000000001100000000000000000000000000000000000100000000000100000000000000100100000000000001010100000000000000000000000000000000000000000001000000000000000100000000000000") port map( O =>C_73_S_0_L_1_out, I0 =>  inp_feat(479), I1 =>  inp_feat(509), I2 =>  inp_feat(234), I3 =>  inp_feat(219), I4 =>  inp_feat(248), I5 =>  inp_feat(68), I6 =>  inp_feat(67), I7 =>  inp_feat(505)); 
C_73_S_0_L_2_inst : LUT8 generic map(INIT => "1111000000000000001000000000000000110000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_0_L_2_out, I0 =>  inp_feat(281), I1 =>  inp_feat(265), I2 =>  inp_feat(400), I3 =>  inp_feat(492), I4 =>  inp_feat(460), I5 =>  inp_feat(240), I6 =>  inp_feat(494), I7 =>  inp_feat(422)); 
C_73_S_0_L_3_inst : LUT8 generic map(INIT => "0001110000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_0_L_3_out, I0 =>  inp_feat(311), I1 =>  inp_feat(72), I2 =>  inp_feat(455), I3 =>  inp_feat(53), I4 =>  inp_feat(504), I5 =>  inp_feat(160), I6 =>  inp_feat(412), I7 =>  inp_feat(58)); 
C_73_S_0_L_4_inst : LUT8 generic map(INIT => "0000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000110000000001010000000000000000000000000001100001000000000000000000111010011001100000000000000100000000010000000000000000000000010000000000110110000000000000000") port map( O =>C_73_S_0_L_4_out, I0 =>  inp_feat(243), I1 =>  inp_feat(381), I2 =>  inp_feat(469), I3 =>  inp_feat(160), I4 =>  inp_feat(303), I5 =>  inp_feat(323), I6 =>  inp_feat(437), I7 =>  inp_feat(167)); 
C_73_S_0_L_5_inst : LUT8 generic map(INIT => "0100001000000010000001000000001010100110000000000000000000000000000000000000001000100000000000001010001000000000000000000000000000100010001000100010000000100000001000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000") port map( O =>C_73_S_0_L_5_out, I0 =>  inp_feat(161), I1 =>  inp_feat(461), I2 =>  inp_feat(437), I3 =>  inp_feat(398), I4 =>  inp_feat(501), I5 =>  inp_feat(348), I6 =>  inp_feat(107), I7 =>  inp_feat(434)); 
C_73_S_0_L_6_inst : LUT8 generic map(INIT => "1010101100000000100010110000000000000000000000000010001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_0_L_6_out, I0 =>  inp_feat(16), I1 =>  inp_feat(483), I2 =>  inp_feat(469), I3 =>  inp_feat(494), I4 =>  inp_feat(308), I5 =>  inp_feat(166), I6 =>  inp_feat(412), I7 =>  inp_feat(240)); 
C_73_S_0_L_7_inst : LUT8 generic map(INIT => "1111001100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011000000001100000000000000010000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_0_L_7_out, I0 =>  inp_feat(437), I1 =>  inp_feat(338), I2 =>  inp_feat(434), I3 =>  inp_feat(128), I4 =>  inp_feat(388), I5 =>  inp_feat(58), I6 =>  inp_feat(420), I7 =>  inp_feat(80)); 
C_73_S_1_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000001000001000000000000000000000000000000000001000000000000000000000000010100000000000001010000000000000101000000000000000100000000000001010000000000000") port map( O =>C_73_S_1_L_0_out, I0 =>  inp_feat(128), I1 =>  inp_feat(351), I2 =>  inp_feat(178), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_73_S_1_L_1_inst : LUT8 generic map(INIT => "0000000000001000000000000000000000001000000010000000100010001000000000000000000000000000000000000000100010000000000000000000000000000000000010001000100000000000000000001000000000001000100010000000000000000000000000000000000000001000000000001000100000000000") port map( O =>C_73_S_1_L_1_out, I0 =>  inp_feat(98), I1 =>  inp_feat(123), I2 =>  inp_feat(237), I3 =>  inp_feat(186), I4 =>  inp_feat(248), I5 =>  inp_feat(68), I6 =>  inp_feat(67), I7 =>  inp_feat(505)); 
C_73_S_1_L_2_inst : LUT8 generic map(INIT => "1100110010100100101010000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_1_L_2_out, I0 =>  inp_feat(394), I1 =>  inp_feat(332), I2 =>  inp_feat(382), I3 =>  inp_feat(437), I4 =>  inp_feat(241), I5 =>  inp_feat(494), I6 =>  inp_feat(219), I7 =>  inp_feat(422)); 
C_73_S_1_L_3_inst : LUT8 generic map(INIT => "0110100000000010110010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_1_L_3_out, I0 =>  inp_feat(303), I1 =>  inp_feat(363), I2 =>  inp_feat(234), I3 =>  inp_feat(58), I4 =>  inp_feat(381), I5 =>  inp_feat(232), I6 =>  inp_feat(412), I7 =>  inp_feat(492)); 
C_73_S_1_L_4_inst : LUT8 generic map(INIT => "0000001000001110000000000000000010110011111000100000000000000000000000000000000000000111000000000000000000000010000000000000000010001010100000000000000000000000001100111010001000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_1_L_4_out, I0 =>  inp_feat(340), I1 =>  inp_feat(343), I2 =>  inp_feat(364), I3 =>  inp_feat(437), I4 =>  inp_feat(128), I5 =>  inp_feat(80), I6 =>  inp_feat(501), I7 =>  inp_feat(348)); 
C_73_S_1_L_5_inst : LUT8 generic map(INIT => "0000000000000011000001100101001100000000000000000000000000000000000100000111000100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000010000000000000100000000000000000000000000000000") port map( O =>C_73_S_1_L_5_out, I0 =>  inp_feat(190), I1 =>  inp_feat(351), I2 =>  inp_feat(206), I3 =>  inp_feat(281), I4 =>  inp_feat(6), I5 =>  inp_feat(57), I6 =>  inp_feat(505), I7 =>  inp_feat(22)); 
C_73_S_1_L_6_inst : LUT8 generic map(INIT => "1100000000000000100000000000000000000000000000001100000000000000100000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_1_L_6_out, I0 =>  inp_feat(115), I1 =>  inp_feat(400), I2 =>  inp_feat(123), I3 =>  inp_feat(504), I4 =>  inp_feat(237), I5 =>  inp_feat(245), I6 =>  inp_feat(437), I7 =>  inp_feat(412)); 
C_73_S_1_L_7_inst : LUT8 generic map(INIT => "0010001010001000101010100000101000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_1_L_7_out, I0 =>  inp_feat(504), I1 =>  inp_feat(281), I2 =>  inp_feat(338), I3 =>  inp_feat(223), I4 =>  inp_feat(505), I5 =>  inp_feat(494), I6 =>  inp_feat(198), I7 =>  inp_feat(422)); 
C_73_S_2_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000001000001000000000000000000000000000000000001000000000000000000000000010100000000000001010000000000000101000000000000000100000000000001010000000000000") port map( O =>C_73_S_2_L_0_out, I0 =>  inp_feat(128), I1 =>  inp_feat(351), I2 =>  inp_feat(178), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_73_S_2_L_1_inst : LUT8 generic map(INIT => "1100110010001100000000000000000000000000000010000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_1_out, I0 =>  inp_feat(432), I1 =>  inp_feat(504), I2 =>  inp_feat(206), I3 =>  inp_feat(308), I4 =>  inp_feat(492), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_73_S_2_L_2_inst : LUT8 generic map(INIT => "0000010100000001000100010000000100000000000000000000100101010001000000000000000000000000000000000000000000000000000000000000000000000011000000000100000000010001000000000001100000010000000100010000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_2_out, I0 =>  inp_feat(281), I1 =>  inp_feat(167), I2 =>  inp_feat(505), I3 =>  inp_feat(348), I4 =>  inp_feat(381), I5 =>  inp_feat(243), I6 =>  inp_feat(422), I7 =>  inp_feat(43)); 
C_73_S_2_L_3_inst : LUT8 generic map(INIT => "0010000000101010000000000000000000000000000000000000000000000000101000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(406), I2 =>  inp_feat(85), I3 =>  inp_feat(243), I4 =>  inp_feat(219), I5 =>  inp_feat(422), I6 =>  inp_feat(43), I7 =>  inp_feat(481)); 
C_73_S_2_L_4_inst : LUT8 generic map(INIT => "0010001000101000101000100000000000100000100000001010000000100000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_4_out, I0 =>  inp_feat(504), I1 =>  inp_feat(80), I2 =>  inp_feat(383), I3 =>  inp_feat(350), I4 =>  inp_feat(381), I5 =>  inp_feat(243), I6 =>  inp_feat(470), I7 =>  inp_feat(313)); 
C_73_S_2_L_5_inst : LUT8 generic map(INIT => "0000100000001000100010000000100000000000000000001000000010100000000000100000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_5_out, I0 =>  inp_feat(494), I1 =>  inp_feat(303), I2 =>  inp_feat(479), I3 =>  inp_feat(346), I4 =>  inp_feat(308), I5 =>  inp_feat(75), I6 =>  inp_feat(313), I7 =>  inp_feat(460)); 
C_73_S_2_L_6_inst : LUT8 generic map(INIT => "0000000000101010101010001000101010001000001010100000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_6_out, I0 =>  inp_feat(494), I1 =>  inp_feat(353), I2 =>  inp_feat(237), I3 =>  inp_feat(406), I4 =>  inp_feat(339), I5 =>  inp_feat(408), I6 =>  inp_feat(422), I7 =>  inp_feat(460)); 
C_73_S_2_L_7_inst : LUT8 generic map(INIT => "0110000000000000000000000010000000010000000000000010000000100000000000000000000000001000101000000000000000001000000000000010000000000000101000001010000000100000000000000000000000100000001000000000000000000000001000000000000000000000000000000000000000000000") port map( O =>C_73_S_2_L_7_out, I0 =>  inp_feat(388), I1 =>  inp_feat(80), I2 =>  inp_feat(312), I3 =>  inp_feat(327), I4 =>  inp_feat(265), I5 =>  inp_feat(508), I6 =>  inp_feat(280), I7 =>  inp_feat(372)); 
C_73_S_3_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000001000001000000000000000000000000000000000001000000000000000000000000010100000000000001010000000000000101000000000000000100000000000001010000000000000") port map( O =>C_73_S_3_L_0_out, I0 =>  inp_feat(128), I1 =>  inp_feat(351), I2 =>  inp_feat(178), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_73_S_3_L_1_inst : LUT8 generic map(INIT => "1100110010001100000000000000000000000000000010000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_3_L_1_out, I0 =>  inp_feat(432), I1 =>  inp_feat(504), I2 =>  inp_feat(206), I3 =>  inp_feat(308), I4 =>  inp_feat(492), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_73_S_3_L_2_inst : LUT8 generic map(INIT => "0001010100000000000100110000000000000000000000001111100100000000000000000000000000000000000000000000000000000000000000000000000001010000000000000001100100000000000100010000000011110000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_3_L_2_out, I0 =>  inp_feat(338), I1 =>  inp_feat(406), I2 =>  inp_feat(437), I3 =>  inp_feat(276), I4 =>  inp_feat(381), I5 =>  inp_feat(243), I6 =>  inp_feat(422), I7 =>  inp_feat(43)); 
C_73_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000000000100000000000000010001000000000001000100000001000000000000000000000000000000000000000000000000000000000000000000010101000000000000000000000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_3_L_3_out, I0 =>  inp_feat(400), I1 =>  inp_feat(170), I2 =>  inp_feat(437), I3 =>  inp_feat(494), I4 =>  inp_feat(505), I5 =>  inp_feat(455), I6 =>  inp_feat(219), I7 =>  inp_feat(160)); 
C_73_S_3_L_4_inst : LUT8 generic map(INIT => "0000000000001000000000000000000011110001000000000000000000000000101010000000000000000000100000000010001110100010000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_3_L_4_out, I0 =>  inp_feat(434), I1 =>  inp_feat(167), I2 =>  inp_feat(340), I3 =>  inp_feat(508), I4 =>  inp_feat(170), I5 =>  inp_feat(455), I6 =>  inp_feat(160), I7 =>  inp_feat(128)); 
C_73_S_3_L_5_inst : LUT8 generic map(INIT => "0101000010010000110000001101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_3_L_5_out, I0 =>  inp_feat(444), I1 =>  inp_feat(162), I2 =>  inp_feat(494), I3 =>  inp_feat(437), I4 =>  inp_feat(237), I5 =>  inp_feat(128), I6 =>  inp_feat(422), I7 =>  inp_feat(359)); 
C_73_S_3_L_6_inst : LUT8 generic map(INIT => "0011000010100000000000000000000000000000000000000000000000000000000100000010100000100000000000000000000000000000000000000000000010000000101100001010100000110000000000000000000000000000000000000000000010100000000000000010000000000000000000000000000000000000") port map( O =>C_73_S_3_L_6_out, I0 =>  inp_feat(434), I1 =>  inp_feat(479), I2 =>  inp_feat(232), I3 =>  inp_feat(237), I4 =>  inp_feat(107), I5 =>  inp_feat(422), I6 =>  inp_feat(359), I7 =>  inp_feat(190)); 
C_73_S_3_L_7_inst : LUT8 generic map(INIT => "0110000000001100000000001000000000000000100001110000000000000100100111001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_3_L_7_out, I0 =>  inp_feat(483), I1 =>  inp_feat(176), I2 =>  inp_feat(478), I3 =>  inp_feat(265), I4 =>  inp_feat(460), I5 =>  inp_feat(128), I6 =>  inp_feat(459), I7 =>  inp_feat(503)); 
C_73_S_4_L_0_inst : LUT8 generic map(INIT => "0000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000001000001000000000000000000000000000000000001000000000000000000000000010100000000000001010000000000000101000000000000000100000000000001010000000000000") port map( O =>C_73_S_4_L_0_out, I0 =>  inp_feat(128), I1 =>  inp_feat(351), I2 =>  inp_feat(178), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_73_S_4_L_1_inst : LUT8 generic map(INIT => "1110000010000000101000001010000000000000000000000000000010000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_4_L_1_out, I0 =>  inp_feat(128), I1 =>  inp_feat(339), I2 =>  inp_feat(504), I3 =>  inp_feat(206), I4 =>  inp_feat(308), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_73_S_4_L_2_inst : LUT8 generic map(INIT => "0001000100000000000000000000000000010001000000001101010100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010010000000000000110010000000011010000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_4_L_2_out, I0 =>  inp_feat(194), I1 =>  inp_feat(336), I2 =>  inp_feat(437), I3 =>  inp_feat(276), I4 =>  inp_feat(243), I5 =>  inp_feat(381), I6 =>  inp_feat(422), I7 =>  inp_feat(43)); 
C_73_S_4_L_3_inst : LUT8 generic map(INIT => "0000000010000000000000001000100010000000100000000000000000000000100000001000100000000000000000001000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_4_L_3_out, I0 =>  inp_feat(422), I1 =>  inp_feat(412), I2 =>  inp_feat(88), I3 =>  inp_feat(413), I4 =>  inp_feat(240), I5 =>  inp_feat(348), I6 =>  inp_feat(483), I7 =>  inp_feat(492)); 
C_73_S_4_L_4_inst : LUT8 generic map(INIT => "0000000000000000000000000110000000000000000000000000000000000000000000000100000010000000110100000000000000000000000000000000000011000000110000000100000001000000000000000000000000000000000000001100000001000000010000000100000000000000000000000000000000000000") port map( O =>C_73_S_4_L_4_out, I0 =>  inp_feat(167), I1 =>  inp_feat(460), I2 =>  inp_feat(412), I3 =>  inp_feat(505), I4 =>  inp_feat(467), I5 =>  inp_feat(400), I6 =>  inp_feat(220), I7 =>  inp_feat(381)); 
C_73_S_4_L_5_inst : LUT8 generic map(INIT => "0000000000000000000010000000000000000000000000000010101000000000100010000000000010001000000000000000000000000000000000000000000010000000000010001000100000000000000000000000000000000000000000000000100000000000100010000000000000000000000000000000000000000000") port map( O =>C_73_S_4_L_5_out, I0 =>  inp_feat(235), I1 =>  inp_feat(141), I2 =>  inp_feat(206), I3 =>  inp_feat(494), I4 =>  inp_feat(351), I5 =>  inp_feat(27), I6 =>  inp_feat(473), I7 =>  inp_feat(505)); 
C_73_S_4_L_6_inst : LUT8 generic map(INIT => "0000000000000010100001101000101000000000000000001000000010001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_73_S_4_L_6_out, I0 =>  inp_feat(494), I1 =>  inp_feat(131), I2 =>  inp_feat(467), I3 =>  inp_feat(167), I4 =>  inp_feat(281), I5 =>  inp_feat(499), I6 =>  inp_feat(198), I7 =>  inp_feat(378)); 
C_73_S_4_L_7_inst : LUT8 generic map(INIT => "0110000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000010000000000000000000000010000001100000000000000000000000000000000000000000000000000000000000000001000000000000000000000") port map( O =>C_73_S_4_L_7_out, I0 =>  inp_feat(167), I1 =>  inp_feat(337), I2 =>  inp_feat(345), I3 =>  inp_feat(280), I4 =>  inp_feat(422), I5 =>  inp_feat(297), I6 =>  inp_feat(494), I7 =>  inp_feat(339)); 
C_74_S_0_L_0_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_1_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_2_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_3_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_4_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_5_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_6_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_0_L_7_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_0_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_0_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_1_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_2_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_3_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_4_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_5_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_6_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_1_L_7_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_1_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_0_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_1_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_2_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_3_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_4_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_5_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_6_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_2_L_7_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_2_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_0_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_1_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_2_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_3_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_4_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_5_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_6_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_3_L_7_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_3_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_0_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_1_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_2_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_3_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_4_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_5_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_6_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_6_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_74_S_4_L_7_inst : LUT8 generic map(INIT => "1111100011100000111010000000100011111000000000001111101000000000111000001110000000000000000000001110000001010000000000000000000011000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_74_S_4_L_7_out, I0 =>  inp_feat(1), I1 =>  inp_feat(0), I2 =>  inp_feat(22), I3 =>  inp_feat(473), I4 =>  inp_feat(68), I5 =>  inp_feat(180), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_75_S_0_L_0_inst : LUT8 generic map(INIT => "1111111011000000101011101010000011110000100100001010000000000000111010001100000010100000111000000000000000000000000000000000000010101010001000001010000010100000101000100000000010100000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_0_L_0_out, I0 =>  inp_feat(241), I1 =>  inp_feat(375), I2 =>  inp_feat(132), I3 =>  inp_feat(80), I4 =>  inp_feat(366), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_75_S_0_L_1_inst : LUT8 generic map(INIT => "0010000000100010111000001000000011100000001000101100000000000000111001001011000010000000000000001111000000000000000000000000000011101000001000101110000010000000111000001110101011000000110000001111111101110101000000000000000010110000000000000000000000000000") port map( O =>C_75_S_0_L_1_out, I0 =>  inp_feat(206), I1 =>  inp_feat(475), I2 =>  inp_feat(339), I3 =>  inp_feat(153), I4 =>  inp_feat(240), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_75_S_0_L_2_inst : LUT8 generic map(INIT => "1111101010101010111110101010101000001000100000001000100010000000100010001000000010001000000000001000100010000000000010000000000000001000101010000000100010000000000000001000000000000000100000001000100000000000000010000000000000001000000000000000100000000000") port map( O =>C_75_S_0_L_2_out, I0 =>  inp_feat(206), I1 =>  inp_feat(237), I2 =>  inp_feat(223), I3 =>  inp_feat(400), I4 =>  inp_feat(379), I5 =>  inp_feat(505), I6 =>  inp_feat(219), I7 =>  inp_feat(455)); 
C_75_S_0_L_3_inst : LUT8 generic map(INIT => "1011111110001011101010001000000011001000000011001000100000001100111111110001000110100000000000001000000000000000100000001000000010001111000001101001110000000000100010000000110000001000000011001111111100000001101000000000000010000000000000000000000000000000") port map( O =>C_75_S_0_L_3_out, I0 =>  inp_feat(281), I1 =>  inp_feat(331), I2 =>  inp_feat(27), I3 =>  inp_feat(357), I4 =>  inp_feat(221), I5 =>  inp_feat(434), I6 =>  inp_feat(120), I7 =>  inp_feat(483)); 
C_75_S_0_L_4_inst : LUT8 generic map(INIT => "1111011111110111111111011101111111000000110100000100000000000000011101010111000000000000000000001100000001000000000000000000000010110011001100110000000000011011000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_0_L_4_out, I0 =>  inp_feat(494), I1 =>  inp_feat(221), I2 =>  inp_feat(467), I3 =>  inp_feat(121), I4 =>  inp_feat(43), I5 =>  inp_feat(381), I6 =>  inp_feat(206), I7 =>  inp_feat(243)); 
C_75_S_0_L_5_inst : LUT8 generic map(INIT => "1101110011001100111111000000110000001100000010001000111100001111110010001000100000000000000010000000000000001000000000000000000000000000000010000000100000001000000000000000100000001000000010001000000010001000000000001000100000000000100010000000000000001000") port map( O =>C_75_S_0_L_5_out, I0 =>  inp_feat(504), I1 =>  inp_feat(80), I2 =>  inp_feat(329), I3 =>  inp_feat(221), I4 =>  inp_feat(128), I5 =>  inp_feat(114), I6 =>  inp_feat(486), I7 =>  inp_feat(243)); 
C_75_S_0_L_6_inst : LUT8 generic map(INIT => "1011100011111000111110101110010000101000111100001111000000100000000000000100000011100010101100000000000000000100110101010101011110001000100010001000100010000000000010001000100010001000100010001000100011000100100000001100001000000100010011001100001011010101") port map( O =>C_75_S_0_L_6_out, I0 =>  inp_feat(281), I1 =>  inp_feat(93), I2 =>  inp_feat(280), I3 =>  inp_feat(504), I4 =>  inp_feat(494), I5 =>  inp_feat(80), I6 =>  inp_feat(155), I7 =>  inp_feat(375)); 
C_75_S_0_L_7_inst : LUT8 generic map(INIT => "0100111010001001110010000000000011101111101001000000000000000000110010000010100000001000000000000000000000000000000000000000000011001101101111011100100010001000111011011110010100000000000000000000100010001000110010000000000000000000000000000000000000000000") port map( O =>C_75_S_0_L_7_out, I0 =>  inp_feat(80), I1 =>  inp_feat(337), I2 =>  inp_feat(494), I3 =>  inp_feat(357), I4 =>  inp_feat(398), I5 =>  inp_feat(375), I6 =>  inp_feat(505), I7 =>  inp_feat(232)); 
C_75_S_1_L_0_inst : LUT8 generic map(INIT => "1111111011000000101011101010000011110000100100001010000000000000111010001100000010100000111000000000000000000000000000000000000010101010001000001010000010100000101000100000000010100000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_1_L_0_out, I0 =>  inp_feat(241), I1 =>  inp_feat(375), I2 =>  inp_feat(132), I3 =>  inp_feat(80), I4 =>  inp_feat(366), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_75_S_1_L_1_inst : LUT8 generic map(INIT => "0010000000100010111000001000000011100000001000101100000000000000111001001011000010000000000000001111000000000000000000000000000011101000001000101110000010000000111000001110101011000000110000001111111101110101000000000000000010110000000000000000000000000000") port map( O =>C_75_S_1_L_1_out, I0 =>  inp_feat(206), I1 =>  inp_feat(475), I2 =>  inp_feat(339), I3 =>  inp_feat(153), I4 =>  inp_feat(240), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_75_S_1_L_2_inst : LUT8 generic map(INIT => "1111101010101010111110101010101000001000100000001000100010000000100010001000000010001000000000001000100010000000000010000000000000001000101010000000100010000000000000001000000000000000100000001000100000000000000010000000000000001000000000000000100000000000") port map( O =>C_75_S_1_L_2_out, I0 =>  inp_feat(206), I1 =>  inp_feat(237), I2 =>  inp_feat(223), I3 =>  inp_feat(400), I4 =>  inp_feat(379), I5 =>  inp_feat(505), I6 =>  inp_feat(219), I7 =>  inp_feat(455)); 
C_75_S_1_L_3_inst : LUT8 generic map(INIT => "1111110111011001111010100000100000000000000000001000001000001000111101111110101010101010101010101111000010100000100000001000101000000000000000000000000000000000000000000000000000000000000000001010000010000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_1_L_3_out, I0 =>  inp_feat(350), I1 =>  inp_feat(379), I2 =>  inp_feat(461), I3 =>  inp_feat(356), I4 =>  inp_feat(400), I5 =>  inp_feat(455), I6 =>  inp_feat(494), I7 =>  inp_feat(160)); 
C_75_S_1_L_4_inst : LUT8 generic map(INIT => "1111111011100110111100111111011110100000001100001000000000000000011010101011001011110101001100110011000011110000111100000111001010001110100000000000001000000010000000000000000000000000000000001000101000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_1_L_4_out, I0 =>  inp_feat(375), I1 =>  inp_feat(494), I2 =>  inp_feat(221), I3 =>  inp_feat(483), I4 =>  inp_feat(437), I5 =>  inp_feat(381), I6 =>  inp_feat(413), I7 =>  inp_feat(243)); 
C_75_S_1_L_5_inst : LUT8 generic map(INIT => "1101110010111100010000001111100010001000000010000010000010001000111010000000100000000000000000000000000000000000000000000000000000011000000000000000000000000000101010000000000010010000000000001111100000000000010000000000000011110000000000001110000000000000") port map( O =>C_75_S_1_L_5_out, I0 =>  inp_feat(274), I1 =>  inp_feat(25), I2 =>  inp_feat(58), I3 =>  inp_feat(20), I4 =>  inp_feat(234), I5 =>  inp_feat(375), I6 =>  inp_feat(422), I7 =>  inp_feat(508)); 
C_75_S_1_L_6_inst : LUT8 generic map(INIT => "0110111010101110010001001100110010101010101010100100000011000000000000001000100000000000000000001010100000101010000000000000000011100100111000000000000010000000110000001100000001000000110000000000000000000000000000000000000000100000110000000000000000000000") port map( O =>C_75_S_1_L_6_out, I0 =>  inp_feat(486), I1 =>  inp_feat(480), I2 =>  inp_feat(169), I3 =>  inp_feat(228), I4 =>  inp_feat(25), I5 =>  inp_feat(375), I6 =>  inp_feat(206), I7 =>  inp_feat(422)); 
C_75_S_1_L_7_inst : LUT8 generic map(INIT => "1111110011110100111101001110110011001000100000001100000010000000000000001111000011000000110000000000000010000000100000001000000001101000110000000000000010000000100000001000000010000000100000001000000010000000000000000000000010000000100000000000000010000000") port map( O =>C_75_S_1_L_7_out, I0 =>  inp_feat(238), I1 =>  inp_feat(80), I2 =>  inp_feat(234), I3 =>  inp_feat(176), I4 =>  inp_feat(166), I5 =>  inp_feat(191), I6 =>  inp_feat(505), I7 =>  inp_feat(23)); 
C_75_S_2_L_0_inst : LUT8 generic map(INIT => "1111111011000000101011101010000011110000100100001010000000000000111010001100000010100000111000000000000000000000000000000000000010101010001000001010000010100000101000100000000010100000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_2_L_0_out, I0 =>  inp_feat(241), I1 =>  inp_feat(375), I2 =>  inp_feat(132), I3 =>  inp_feat(80), I4 =>  inp_feat(366), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_75_S_2_L_1_inst : LUT8 generic map(INIT => "0010000000100010111000001000000011100000001000101100000000000000111001001011000010000000000000001111000000000000000000000000000011101000001000101110000010000000111000001110101011000000110000001111111101110101000000000000000010110000000000000000000000000000") port map( O =>C_75_S_2_L_1_out, I0 =>  inp_feat(206), I1 =>  inp_feat(475), I2 =>  inp_feat(339), I3 =>  inp_feat(153), I4 =>  inp_feat(240), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_75_S_2_L_2_inst : LUT8 generic map(INIT => "1111011011111100101110111101100110001010111110001011111111011010101100000011000010001111000000001000000001110000101101011000100010100000100000001010100010001000101000100000000010100001000000000000000000000000000011000000100000000000000000001010000000000000") port map( O =>C_75_S_2_L_2_out, I0 =>  inp_feat(479), I1 =>  inp_feat(379), I2 =>  inp_feat(6), I3 =>  inp_feat(474), I4 =>  inp_feat(72), I5 =>  inp_feat(166), I6 =>  inp_feat(505), I7 =>  inp_feat(455)); 
C_75_S_2_L_3_inst : LUT8 generic map(INIT => "1000100110110000111101101111000010101100101000001110111001000000000000000010000001000000000000001010000010100000110000000100000010000000100000001100000011000000101000101000000010100000000000000000000010000000010000000000000000000000100000000000000000000000") port map( O =>C_75_S_2_L_3_out, I0 =>  inp_feat(408), I1 =>  inp_feat(149), I2 =>  inp_feat(206), I3 =>  inp_feat(311), I4 =>  inp_feat(232), I5 =>  inp_feat(399), I6 =>  inp_feat(243), I7 =>  inp_feat(486)); 
C_75_S_2_L_4_inst : LUT8 generic map(INIT => "1110111011001100111011101100101001101110110010001110111100000010110011001100110010000010100010100000000000000000000010100000101011000000110001000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_2_L_4_out, I0 =>  inp_feat(340), I1 =>  inp_feat(508), I2 =>  inp_feat(102), I3 =>  inp_feat(494), I4 =>  inp_feat(332), I5 =>  inp_feat(68), I6 =>  inp_feat(80), I7 =>  inp_feat(451)); 
C_75_S_2_L_5_inst : LUT8 generic map(INIT => "1000110001001110111100000000000010000100000011000001000000000000111111111111111111010011001100110111110000011100100100000000000011001100100011001100000000000000000011000000101000000000000000001000000010010000100000000000000000000000100000000000000000000000") port map( O =>C_75_S_2_L_5_out, I0 =>  inp_feat(290), I1 =>  inp_feat(281), I2 =>  inp_feat(58), I3 =>  inp_feat(238), I4 =>  inp_feat(357), I5 =>  inp_feat(206), I6 =>  inp_feat(102), I7 =>  inp_feat(221)); 
C_75_S_2_L_6_inst : LUT8 generic map(INIT => "1111011110100000101010101010000001010000101000001010000010100000111111111010001110000000101000000010000010100000101000001010000000110011100000001000100010000000000000001000000000000000000000001011001111110011100000001000000010000000110000001000000010000000") port map( O =>C_75_S_2_L_6_out, I0 =>  inp_feat(503), I1 =>  inp_feat(375), I2 =>  inp_feat(234), I3 =>  inp_feat(504), I4 =>  inp_feat(494), I5 =>  inp_feat(80), I6 =>  inp_feat(379), I7 =>  inp_feat(34)); 
C_75_S_2_L_7_inst : LUT8 generic map(INIT => "1010001011000000111010101100000011110010000000001010001010000000111100001000000010010000110000001000000010000000000000001000000011111011110000011111101111001111111100001000000010000000100000001010000011100000000000001100000010100000001000001000000010000000") port map( O =>C_75_S_2_L_7_out, I0 =>  inp_feat(190), I1 =>  inp_feat(385), I2 =>  inp_feat(237), I3 =>  inp_feat(19), I4 =>  inp_feat(379), I5 =>  inp_feat(351), I6 =>  inp_feat(166), I7 =>  inp_feat(176)); 
C_75_S_3_L_0_inst : LUT8 generic map(INIT => "1111111011000000101011101010000011110000100100001010000000000000111010001100000010100000111000000000000000000000000000000000000010101010001000001010000010100000101000100000000010100000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_3_L_0_out, I0 =>  inp_feat(241), I1 =>  inp_feat(375), I2 =>  inp_feat(132), I3 =>  inp_feat(80), I4 =>  inp_feat(366), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_75_S_3_L_1_inst : LUT8 generic map(INIT => "0010000000100010111000001000000011100000001000101100000000000000111001001011000010000000000000001111000000000000000000000000000011101000001000101110000010000000111000001110101011000000110000001111111101110101000000000000000010110000000000000000000000000000") port map( O =>C_75_S_3_L_1_out, I0 =>  inp_feat(206), I1 =>  inp_feat(475), I2 =>  inp_feat(339), I3 =>  inp_feat(153), I4 =>  inp_feat(240), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_75_S_3_L_2_inst : LUT8 generic map(INIT => "1111011011111100101110111101100110001010111110001011111111011010101100000011000010001111000000001000000001110000101101011000100010100000100000001010100010001000101000100000000010100001000000000000000000000000000011000000100000000000000000001010000000000000") port map( O =>C_75_S_3_L_2_out, I0 =>  inp_feat(479), I1 =>  inp_feat(379), I2 =>  inp_feat(6), I3 =>  inp_feat(474), I4 =>  inp_feat(72), I5 =>  inp_feat(166), I6 =>  inp_feat(505), I7 =>  inp_feat(455)); 
C_75_S_3_L_3_inst : LUT8 generic map(INIT => "1011110010000000111011101000100010100000100000001000100010000000100001000000000010001000000000001010000000000000100000000000000011100000100000001000100010000000101000000000000010000000100000000010000000000000100000001000000010100000000000001000000000000000") port map( O =>C_75_S_3_L_3_out, I0 =>  inp_feat(206), I1 =>  inp_feat(180), I2 =>  inp_feat(483), I3 =>  inp_feat(381), I4 =>  inp_feat(232), I5 =>  inp_feat(219), I6 =>  inp_feat(243), I7 =>  inp_feat(486)); 
C_75_S_3_L_4_inst : LUT8 generic map(INIT => "1011110010111110101000001010000010100000101000000000000000000000111000001110000011000000100000000000000010000000100000000000000010000000101000001010000000000000000000001010000000000000000000001010000010100000100000000000000010000000101000001000000000000000") port map( O =>C_75_S_3_L_4_out, I0 =>  inp_feat(237), I1 =>  inp_feat(68), I2 =>  inp_feat(67), I3 =>  inp_feat(303), I4 =>  inp_feat(503), I5 =>  inp_feat(114), I6 =>  inp_feat(399), I7 =>  inp_feat(243)); 
C_75_S_3_L_5_inst : LUT8 generic map(INIT => "0110111000100010111111000111000001000100000000100000110000000000111111101010101001111111111100000000001010101110001111110101101111101110101010101100110001001000000001000000000011000100000000000000101000000010000000000000000000000000000000000000101000001000") port map( O =>C_75_S_3_L_5_out, I0 =>  inp_feat(375), I1 =>  inp_feat(232), I2 =>  inp_feat(494), I3 =>  inp_feat(265), I4 =>  inp_feat(65), I5 =>  inp_feat(80), I6 =>  inp_feat(102), I7 =>  inp_feat(221)); 
C_75_S_3_L_6_inst : LUT8 generic map(INIT => "1101011111001111110010001100100001000000010000001100110001001100111111111100111111001100010011001100000001000000000000000100000011011110100011100000110000001100110001000100010001000100000011001111111100001100000000000000000011001000000001001100000000000000") port map( O =>C_75_S_3_L_6_out, I0 =>  inp_feat(494), I1 =>  inp_feat(505), I2 =>  inp_feat(468), I3 =>  inp_feat(141), I4 =>  inp_feat(375), I5 =>  inp_feat(206), I6 =>  inp_feat(379), I7 =>  inp_feat(88)); 
C_75_S_3_L_7_inst : LUT8 generic map(INIT => "1111101110110011101000100010000000100000111100000000000000000000001000101010000010100000001000000000000000100000001000000010000011101011000000001000000000000000110000000000000010000000000000001010000010000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_3_L_7_out, I0 =>  inp_feat(25), I1 =>  inp_feat(494), I2 =>  inp_feat(129), I3 =>  inp_feat(20), I4 =>  inp_feat(206), I5 =>  inp_feat(234), I6 =>  inp_feat(374), I7 =>  inp_feat(422)); 
C_75_S_4_L_0_inst : LUT8 generic map(INIT => "1111111011000000101011101010000011110000100100001010000000000000111010001100000010100000111000000000000000000000000000000000000010101010001000001010000010100000101000100000000010100000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_4_L_0_out, I0 =>  inp_feat(241), I1 =>  inp_feat(375), I2 =>  inp_feat(132), I3 =>  inp_feat(80), I4 =>  inp_feat(366), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_75_S_4_L_1_inst : LUT8 generic map(INIT => "0010111100100000000000100010000010101111101010100000000000000011111011001010100010000010000000001010111010101010000010000010100011001101111000011000000100110000110011111000110100000011000001111100000001000000110000000000000011001100000000001000000000000000") port map( O =>C_75_S_4_L_1_out, I0 =>  inp_feat(308), I1 =>  inp_feat(45), I2 =>  inp_feat(217), I3 =>  inp_feat(491), I4 =>  inp_feat(206), I5 =>  inp_feat(98), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_75_S_4_L_2_inst : LUT8 generic map(INIT => "1110111111101100100011001010111010101111001011101010000010101010101010001010101000000000101010001010101000101010101000001010100010100000101000000000000000100000000000000000000000000000000000101000000010100000000000000000000000100000000000000000000000000000") port map( O =>C_75_S_4_L_2_out, I0 =>  inp_feat(206), I1 =>  inp_feat(467), I2 =>  inp_feat(4), I3 =>  inp_feat(379), I4 =>  inp_feat(100), I5 =>  inp_feat(468), I6 =>  inp_feat(505), I7 =>  inp_feat(455)); 
C_75_S_4_L_3_inst : LUT8 generic map(INIT => "0011111110111111101010101010101000100100101001001000000000100000111001001110010000100000101000001010010010100100000000000010000000001110100001001010101000000000000001000000010000000000000000001100010001000000000000000000000000000100000001000000000000000000") port map( O =>C_75_S_4_L_3_out, I0 =>  inp_feat(248), I1 =>  inp_feat(379), I2 =>  inp_feat(240), I3 =>  inp_feat(340), I4 =>  inp_feat(232), I5 =>  inp_feat(243), I6 =>  inp_feat(15), I7 =>  inp_feat(331)); 
C_75_S_4_L_4_inst : LUT8 generic map(INIT => "1101111110101010110101111110001011101010101001001010001000100000111011111000001000000011000000100010000000100000000000100010001000001000000010000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_75_S_4_L_4_out, I0 =>  inp_feat(219), I1 =>  inp_feat(340), I2 =>  inp_feat(467), I3 =>  inp_feat(483), I4 =>  inp_feat(323), I5 =>  inp_feat(372), I6 =>  inp_feat(91), I7 =>  inp_feat(234)); 
C_75_S_4_L_5_inst : LUT8 generic map(INIT => "1110111010001110101011001010000010001100000001001010011010100010110011001100111000000000100000000000000011000100001000101010001000101100000000001110110010000000100000000000000011101110101000101000000000000000000000000000000000000000000000000010001000100010") port map( O =>C_75_S_4_L_5_out, I0 =>  inp_feat(80), I1 =>  inp_feat(68), I2 =>  inp_feat(241), I3 =>  inp_feat(107), I4 =>  inp_feat(221), I5 =>  inp_feat(230), I6 =>  inp_feat(396), I7 =>  inp_feat(65)); 
C_75_S_4_L_6_inst : LUT8 generic map(INIT => "1101110011000000111111011000000000000000100000001100110100000000111100001000000010000000100000001000000010000000100000000000000011110000100000001010000000000000000000000000000000000000000000001101000000000000100000000000000010000000000000001000000000000000") port map( O =>C_75_S_4_L_6_out, I0 =>  inp_feat(375), I1 =>  inp_feat(47), I2 =>  inp_feat(80), I3 =>  inp_feat(142), I4 =>  inp_feat(332), I5 =>  inp_feat(381), I6 =>  inp_feat(400), I7 =>  inp_feat(268)); 
C_75_S_4_L_7_inst : LUT8 generic map(INIT => "1111001011110000001000101111000010101010110010001010101010000000000000001100000000000000101010000000000010000000001000001000000010101010101000001010000010100000000000001000000000100010100000000000000000100000000000001010000000000000000000000000000010000000") port map( O =>C_75_S_4_L_7_out, I0 =>  inp_feat(215), I1 =>  inp_feat(224), I2 =>  inp_feat(80), I3 =>  inp_feat(221), I4 =>  inp_feat(288), I5 =>  inp_feat(241), I6 =>  inp_feat(243), I7 =>  inp_feat(43)); 
C_76_S_0_L_0_inst : LUT8 generic map(INIT => "1111111110100010011111110000000011111110111110000100000000000000111011001100000001001000000000000000000000000000000000000000000011111111001000100101111100000000100010110000001000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_0_L_0_out, I0 =>  inp_feat(475), I1 =>  inp_feat(385), I2 =>  inp_feat(98), I3 =>  inp_feat(80), I4 =>  inp_feat(234), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_76_S_0_L_1_inst : LUT8 generic map(INIT => "1111110100011010011001001000101010100000100000001000000010000000011100000011000000000000000000001110000010000000000000000000000011110101000010000000000000000010101100001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_0_L_1_out, I0 =>  inp_feat(420), I1 =>  inp_feat(431), I2 =>  inp_feat(271), I3 =>  inp_feat(338), I4 =>  inp_feat(238), I5 =>  inp_feat(219), I6 =>  inp_feat(268), I7 =>  inp_feat(505)); 
C_76_S_0_L_2_inst : LUT8 generic map(INIT => "0111110101111110111101010011010101111101000010000010110000001100110111010101100001011101010101001101110100001000110111000000010001111100000000001110000000000000010001000000000000000100000000001100000000000000110001000000000011001000100010000000000000000000") port map( O =>C_76_S_0_L_2_out, I0 =>  inp_feat(494), I1 =>  inp_feat(58), I2 =>  inp_feat(7), I3 =>  inp_feat(281), I4 =>  inp_feat(351), I5 =>  inp_feat(362), I6 =>  inp_feat(388), I7 =>  inp_feat(505)); 
C_76_S_0_L_3_inst : LUT8 generic map(INIT => "1111111111111111010001010110000010100000101100100000000000100000001101110000010001000101000000001010000000000000000000000000000000000100001100000000000000000000101000000011000000000000000000000000000000000000000000000000000010000000000000000000000000000000") port map( O =>C_76_S_0_L_3_out, I0 =>  inp_feat(128), I1 =>  inp_feat(494), I2 =>  inp_feat(468), I3 =>  inp_feat(291), I4 =>  inp_feat(429), I5 =>  inp_feat(250), I6 =>  inp_feat(362), I7 =>  inp_feat(377)); 
C_76_S_0_L_4_inst : LUT8 generic map(INIT => "0001111101100110011001101010001001000110010000100000000000000000011101111111000000000000001000001111110011110010000000000011000011111011110011100100011011001110010001100100011000000110110011101000100011110010000000000000000001100010011100100000000000000010") port map( O =>C_76_S_0_L_4_out, I0 =>  inp_feat(494), I1 =>  inp_feat(422), I2 =>  inp_feat(388), I3 =>  inp_feat(98), I4 =>  inp_feat(347), I5 =>  inp_feat(274), I6 =>  inp_feat(319), I7 =>  inp_feat(475)); 
C_76_S_0_L_5_inst : LUT8 generic map(INIT => "0101111111111010101010101011101010111000101010100000000010101010110011111001011111111111111111110100000101000101000011011111111100100010100010101000001010000010000000100000001000000000100000100000100000001000101010100000000000000000000000000000000000000000") port map( O =>C_76_S_0_L_5_out, I0 =>  inp_feat(446), I1 =>  inp_feat(468), I2 =>  inp_feat(41), I3 =>  inp_feat(170), I4 =>  inp_feat(102), I5 =>  inp_feat(378), I6 =>  inp_feat(93), I7 =>  inp_feat(352)); 
C_76_S_0_L_6_inst : LUT8 generic map(INIT => "1111111110001000110111000000100011001101100010001100100000000000100110111000100000001000000010001100000000000000110000000000000000001100000000000000000000000000111010100000100000011001000000001100100010001000000000001000000001000000000000000000000000000000") port map( O =>C_76_S_0_L_6_out, I0 =>  inp_feat(507), I1 =>  inp_feat(80), I2 =>  inp_feat(494), I3 =>  inp_feat(256), I4 =>  inp_feat(362), I5 =>  inp_feat(363), I6 =>  inp_feat(66), I7 =>  inp_feat(114)); 
C_76_S_0_L_7_inst : LUT8 generic map(INIT => "0010101100001000001110111000000001001010100000000000000000000000010110110000100010111010100000000111101000001010000000000000000011001010100000000100000010000000110000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_0_L_7_out, I0 =>  inp_feat(101), I1 =>  inp_feat(473), I2 =>  inp_feat(497), I3 =>  inp_feat(261), I4 =>  inp_feat(128), I5 =>  inp_feat(486), I6 =>  inp_feat(475), I7 =>  inp_feat(124)); 
C_76_S_1_L_0_inst : LUT8 generic map(INIT => "1110100011101010101000001110100011000000110010001010000010100000111000001010101001000000101000001100000011001000100000001000000000101000011010001010000010100000111001001100110010100000101000001000101010101010000000001010000011001000110011101000000000000000") port map( O =>C_76_S_1_L_0_out, I0 =>  inp_feat(406), I1 =>  inp_feat(80), I2 =>  inp_feat(206), I3 =>  inp_feat(494), I4 =>  inp_feat(93), I5 =>  inp_feat(475), I6 =>  inp_feat(92), I7 =>  inp_feat(362)); 
C_76_S_1_L_1_inst : LUT8 generic map(INIT => "1111000111010001100000001100110011011001110001011000000011000000111101001000000001000100010000001100010001000100010000000100010011000000110000001000000011000000100000000000000010000000000000000000010000000000000000000100000001000000000000000100000000000000") port map( O =>C_76_S_1_L_1_out, I0 =>  inp_feat(102), I1 =>  inp_feat(508), I2 =>  inp_feat(281), I3 =>  inp_feat(11), I4 =>  inp_feat(430), I5 =>  inp_feat(178), I6 =>  inp_feat(343), I7 =>  inp_feat(505)); 
C_76_S_1_L_2_inst : LUT8 generic map(INIT => "0110101010001010101110101111111010110010000011100000100001001110111100001100000011110000111100000111000000000000000000000000000000101010000000000000000000100010000000100000000000000000000000000000000000000000001000000010000000110000000000000000000000000000") port map( O =>C_76_S_1_L_2_out, I0 =>  inp_feat(47), I1 =>  inp_feat(247), I2 =>  inp_feat(494), I3 =>  inp_feat(66), I4 =>  inp_feat(232), I5 =>  inp_feat(351), I6 =>  inp_feat(118), I7 =>  inp_feat(114)); 
C_76_S_1_L_3_inst : LUT8 generic map(INIT => "1010101010101010110010001000100011101010101010100000000010100100101010001000000011001100110000001110101010001010100010001100010000000000100000001000000010000000100000001000000000000000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_1_L_3_out, I0 =>  inp_feat(381), I1 =>  inp_feat(378), I2 =>  inp_feat(181), I3 =>  inp_feat(447), I4 =>  inp_feat(250), I5 =>  inp_feat(232), I6 =>  inp_feat(66), I7 =>  inp_feat(377)); 
C_76_S_1_L_4_inst : LUT8 generic map(INIT => "0101000110111010000000001010000010001000101110100000000000000000111100011111010011110000111100001010000011111010000100001111001010100010110000000000000000000000001000100000101000000000000000001001000011010000100000001100000010000000100110000000000000001000") port map( O =>C_76_S_1_L_4_out, I0 =>  inp_feat(51), I1 =>  inp_feat(265), I2 =>  inp_feat(281), I3 =>  inp_feat(494), I4 =>  inp_feat(256), I5 =>  inp_feat(285), I6 =>  inp_feat(448), I7 =>  inp_feat(74)); 
C_76_S_1_L_5_inst : LUT8 generic map(INIT => "0111001100101010000010000000000011011000000000001000000000000000111110110000100001001000000000001011001100000000000000000000000010111011001000001000000000000000101110110000000000000000000000001111101110001000000010000000000011111011000000000000000000000000") port map( O =>C_76_S_1_L_5_out, I0 =>  inp_feat(378), I1 =>  inp_feat(400), I2 =>  inp_feat(494), I3 =>  inp_feat(381), I4 =>  inp_feat(429), I5 =>  inp_feat(269), I6 =>  inp_feat(431), I7 =>  inp_feat(232)); 
C_76_S_1_L_6_inst : LUT8 generic map(INIT => "0111001011101010110110001010100000000000011000101100000010000000101110101010101010001000100000000000000000000000000000001000000000010000101000000011000000100000000000001010100000101000101010101011000000100000000100000000000000000000000000000000000000000000") port map( O =>C_76_S_1_L_6_out, I0 =>  inp_feat(76), I1 =>  inp_feat(98), I2 =>  inp_feat(342), I3 =>  inp_feat(494), I4 =>  inp_feat(30), I5 =>  inp_feat(80), I6 =>  inp_feat(239), I7 =>  inp_feat(502)); 
C_76_S_1_L_7_inst : LUT8 generic map(INIT => "0011100011111000111010000100000011100000111000001110000000000000000010001100100010000000000000001010100010000000101010101000000011110000000000001110000010000000111100000000000011000000000000000000000000000000100000000000000000000000000000001000000000000000") port map( O =>C_76_S_1_L_7_out, I0 =>  inp_feat(406), I1 =>  inp_feat(238), I2 =>  inp_feat(80), I3 =>  inp_feat(248), I4 =>  inp_feat(430), I5 =>  inp_feat(284), I6 =>  inp_feat(343), I7 =>  inp_feat(434)); 
C_76_S_2_L_0_inst : LUT8 generic map(INIT => "1101111110011111000001001000111111111111011011010000100000001000000001000000010100001110000010001100010000011100000000000000000011001110000000000000101000000000000001000000010100000000000000001100111100000101110011101000101000000100000001010000000000000000") port map( O =>C_76_S_2_L_0_out, I0 =>  inp_feat(7), I1 =>  inp_feat(469), I2 =>  inp_feat(494), I3 =>  inp_feat(5), I4 =>  inp_feat(80), I5 =>  inp_feat(239), I6 =>  inp_feat(502), I7 =>  inp_feat(250)); 
C_76_S_2_L_1_inst : LUT8 generic map(INIT => "1111001001000000101010001000000011010001100000001000000000000000111110001010000011101000101000001000000000000000100000001000000010111011001000001000000000000000111111110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_2_L_1_out, I0 =>  inp_feat(80), I1 =>  inp_feat(192), I2 =>  inp_feat(238), I3 =>  inp_feat(190), I4 =>  inp_feat(239), I5 =>  inp_feat(502), I6 =>  inp_feat(382), I7 =>  inp_feat(250)); 
C_76_S_2_L_2_inst : LUT8 generic map(INIT => "1111101010111010001010110110001111100000101010000000000000000000111010001000100011100000100010000100000000000000100000001000000011101010100010000000000010001000000000001000000000000000001000001100000010000000100000001000000000000000000000001010000010000000") port map( O =>C_76_S_2_L_2_out, I0 =>  inp_feat(502), I1 =>  inp_feat(382), I2 =>  inp_feat(166), I3 =>  inp_feat(288), I4 =>  inp_feat(100), I5 =>  inp_feat(67), I6 =>  inp_feat(209), I7 =>  inp_feat(74)); 
C_76_S_2_L_3_inst : LUT8 generic map(INIT => "0110110011001101100110101101110001001000110111001100100001000100111111100101100001111010000100001101000001010000110000000101000011111000110100000111001000010000010010001101100000000000000000001111101001010000101110100000000001010000010000000000000000010000") port map( O =>C_76_S_2_L_3_out, I0 =>  inp_feat(65), I1 =>  inp_feat(406), I2 =>  inp_feat(469), I3 =>  inp_feat(330), I4 =>  inp_feat(158), I5 =>  inp_feat(237), I6 =>  inp_feat(207), I7 =>  inp_feat(473)); 
C_76_S_2_L_4_inst : LUT8 generic map(INIT => "1101100011011000000010001000100011011101110110101000111100001110010111101000100010001000000000001011001100001000100110010000000001001110000000000000000000000000000100000001000000000000000000001000100000000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_2_L_4_out, I0 =>  inp_feat(123), I1 =>  inp_feat(110), I2 =>  inp_feat(232), I3 =>  inp_feat(383), I4 =>  inp_feat(80), I5 =>  inp_feat(209), I6 =>  inp_feat(427), I7 =>  inp_feat(132)); 
C_76_S_2_L_5_inst : LUT8 generic map(INIT => "1011111111110011111011111101000010111000000100001001000000000000110111011101010001000101110000000000100000000000000000000000000000011000111100001110000001010000000000000000000000000000000000001001010001010000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_2_L_5_out, I0 =>  inp_feat(303), I1 =>  inp_feat(365), I2 =>  inp_feat(343), I3 =>  inp_feat(434), I4 =>  inp_feat(238), I5 =>  inp_feat(248), I6 =>  inp_feat(396), I7 =>  inp_feat(319)); 
C_76_S_2_L_6_inst : LUT8 generic map(INIT => "1101110111000000111110000100000011110000110000001111000000000000101100000000000010000000000000000010000000000000001000000000000001100000110010001100000000000000111000000100000001110000010000001000000010001000100000000000000000000000000000001000000000000000") port map( O =>C_76_S_2_L_6_out, I0 =>  inp_feat(365), I1 =>  inp_feat(167), I2 =>  inp_feat(348), I3 =>  inp_feat(455), I4 =>  inp_feat(468), I5 =>  inp_feat(61), I6 =>  inp_feat(76), I7 =>  inp_feat(411)); 
C_76_S_2_L_7_inst : LUT8 generic map(INIT => "1011110010001100110011000000110011101100110011101110110010001100111001100000101011001100000001001010101000001010100000000000000011111010000000101000000000000000100110000000000010000000000000000000101000001000000000000000000010101010000010101010000000000000") port map( O =>C_76_S_2_L_7_out, I0 =>  inp_feat(65), I1 =>  inp_feat(61), I2 =>  inp_feat(303), I3 =>  inp_feat(265), I4 =>  inp_feat(110), I5 =>  inp_feat(170), I6 =>  inp_feat(427), I7 =>  inp_feat(378)); 
C_76_S_3_L_0_inst : LUT8 generic map(INIT => "1110101010111000111010101111001011011110110011101000100000000000000000001011101010001010000000100000001011101110000000100001100010001010101000001010000000000000100000000000000000000000000000001010000010001000101010100000001010000000110011100010001000000000") port map( O =>C_76_S_3_L_0_out, I0 =>  inp_feat(409), I1 =>  inp_feat(505), I2 =>  inp_feat(198), I3 =>  inp_feat(178), I4 =>  inp_feat(434), I5 =>  inp_feat(50), I6 =>  inp_feat(461), I7 =>  inp_feat(273)); 
C_76_S_3_L_1_inst : LUT8 generic map(INIT => "0110110000000000101100001000000000000000100000001000000000000000111010100000001011000000000000001110000000000000000000000000000011101011100010101000000010000000101000001000000010000000100000001100001000000010000000000000000000000000000000000000000000000000") port map( O =>C_76_S_3_L_1_out, I0 =>  inp_feat(238), I1 =>  inp_feat(351), I2 =>  inp_feat(248), I3 =>  inp_feat(503), I4 =>  inp_feat(396), I5 =>  inp_feat(319), I6 =>  inp_feat(230), I7 =>  inp_feat(273)); 
C_76_S_3_L_2_inst : LUT8 generic map(INIT => "0111110011011100101010000000100011001000010110001000100000000000010101110101000010000000000000001010100011000000000000000000000011111110011001001010000000000000100000000000000010000000000000001111011101110000000000001000000011111011011101011010100000000000") port map( O =>C_76_S_3_L_2_out, I0 =>  inp_feat(494), I1 =>  inp_feat(461), I2 =>  inp_feat(398), I3 =>  inp_feat(505), I4 =>  inp_feat(503), I5 =>  inp_feat(396), I6 =>  inp_feat(319), I7 =>  inp_feat(273)); 
C_76_S_3_L_3_inst : LUT8 generic map(INIT => "0101100110011100111011111100011101010000110010000000000001000000100111001000001100011011010111111110000000000000000000010000110110000000110011111010000111011111111100000100000000000000010000011000101111001111000011110100111111110011000010110000101100001111") port map( O =>C_76_S_3_L_3_out, I0 =>  inp_feat(224), I1 =>  inp_feat(374), I2 =>  inp_feat(345), I3 =>  inp_feat(400), I4 =>  inp_feat(166), I5 =>  inp_feat(378), I6 =>  inp_feat(366), I7 =>  inp_feat(492)); 
C_76_S_3_L_4_inst : LUT8 generic map(INIT => "1110000011100000100000001000000000001100101000001010000010100000100100001101000000000000000000001110101011001000000000000000000011100000111100001100000000000000101011111010000000000000000000000110010001000000000000000000000001110011000000000000000000000000") port map( O =>C_76_S_3_L_4_out, I0 =>  inp_feat(74), I1 =>  inp_feat(98), I2 =>  inp_feat(80), I3 =>  inp_feat(239), I4 =>  inp_feat(350), I5 =>  inp_feat(201), I6 =>  inp_feat(206), I7 =>  inp_feat(270)); 
C_76_S_3_L_5_inst : LUT8 generic map(INIT => "1110111010000000111111111000000011101101000000001111111110000101110011011000000011011111110111011111010111000000110111111101110100000110000000001101111100010101000011110000000010001111010011111000000000000000010011110100111100001010000000000100110111001101") port map( O =>C_76_S_3_L_5_out, I0 =>  inp_feat(475), I1 =>  inp_feat(347), I2 =>  inp_feat(363), I3 =>  inp_feat(66), I4 =>  inp_feat(330), I5 =>  inp_feat(420), I6 =>  inp_feat(7), I7 =>  inp_feat(261)); 
C_76_S_3_L_6_inst : LUT8 generic map(INIT => "0000010011110101111011000100000010100100110001001110010001000000010000000000000000000000000000001100010011000000010000000000000000011101111110101010010000000000110001001100000000000000000000001111000011000000000000000000000011000000110000000000000000000000") port map( O =>C_76_S_3_L_6_out, I0 =>  inp_feat(375), I1 =>  inp_feat(80), I2 =>  inp_feat(206), I3 =>  inp_feat(247), I4 =>  inp_feat(271), I5 =>  inp_feat(475), I6 =>  inp_feat(168), I7 =>  inp_feat(431)); 
C_76_S_3_L_7_inst : LUT8 generic map(INIT => "1110111011100010100000001000100010111010101010100000000000100000001000001000000000000000000000101010101000100010000000000000001011101110111000100100001011000000111010101010101000100010101000101010101000100010000000000000000011101000101000100000000000000010") port map( O =>C_76_S_3_L_7_out, I0 =>  inp_feat(206), I1 =>  inp_feat(276), I2 =>  inp_feat(100), I3 =>  inp_feat(471), I4 =>  inp_feat(502), I5 =>  inp_feat(382), I6 =>  inp_feat(378), I7 =>  inp_feat(98)); 
C_76_S_4_L_0_inst : LUT8 generic map(INIT => "1111100010110001110100000000000000100000101100001111000100110000110110001111100100000000000100001101100111111101111100011111010100000000100000001000000000000000100000001100000000000000000000001100000001000000000000000000000000000000000000000000000000000000") port map( O =>C_76_S_4_L_0_out, I0 =>  inp_feat(6), I1 =>  inp_feat(276), I2 =>  inp_feat(502), I3 =>  inp_feat(347), I4 =>  inp_feat(76), I5 =>  inp_feat(446), I6 =>  inp_feat(98), I7 =>  inp_feat(62)); 
C_76_S_4_L_1_inst : LUT8 generic map(INIT => "1101110011111100110011000101111010001100100011000000100000001100100000001110000011000000110011001000100010001100000011000000110011000000110010001100100011001111000000000000110000001000000011100000000011100000000000001110100000001000000001000000100000001100") port map( O =>C_76_S_4_L_1_out, I0 =>  inp_feat(352), I1 =>  inp_feat(281), I2 =>  inp_feat(508), I3 =>  inp_feat(232), I4 =>  inp_feat(431), I5 =>  inp_feat(168), I6 =>  inp_feat(473), I7 =>  inp_feat(66)); 
C_76_S_4_L_2_inst : LUT8 generic map(INIT => "1101000011111100110000001110000011001100111111001000100111110000111100001111000010000000100000001000000010010000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011110000100000000000000000000000000000000000000000000000") port map( O =>C_76_S_4_L_2_out, I0 =>  inp_feat(373), I1 =>  inp_feat(238), I2 =>  inp_feat(461), I3 =>  inp_feat(494), I4 =>  inp_feat(193), I5 =>  inp_feat(161), I6 =>  inp_feat(250), I7 =>  inp_feat(377)); 
C_76_S_4_L_3_inst : LUT8 generic map(INIT => "1111101111111011100000001010001010111010000000000000000000000000100010001111101000001010000010101010101000000000001000000000000000111000000000000000100000001000101110000000000000001000000000001000100000000000000010000000100000000000000000000000100000001000") port map( O =>C_76_S_4_L_3_out, I0 =>  inp_feat(357), I1 =>  inp_feat(11), I2 =>  inp_feat(178), I3 =>  inp_feat(30), I4 =>  inp_feat(248), I5 =>  inp_feat(430), I6 =>  inp_feat(74), I7 =>  inp_feat(378)); 
C_76_S_4_L_4_inst : LUT8 generic map(INIT => "1101101000101011000000001010000010001111101011100000000010000000000010000000000010000000100000001000000010000000100000001000000011000010101010100101000000000000101000001010001010000000100000001000000010000000100000001000000010000000100000001000000010000000") port map( O =>C_76_S_4_L_4_out, I0 =>  inp_feat(74), I1 =>  inp_feat(365), I2 =>  inp_feat(128), I3 =>  inp_feat(309), I4 =>  inp_feat(237), I5 =>  inp_feat(475), I6 =>  inp_feat(168), I7 =>  inp_feat(431)); 
C_76_S_4_L_5_inst : LUT8 generic map(INIT => "1110100010101000111111001110100010001000110000000000110011001100101010011010001011111110111111000000000000000000000000000000000000001000000000001100110010000000010001001000000011000000110001001000110010000001011111001110000000000000000000000000000000000000") port map( O =>C_76_S_4_L_5_out, I0 =>  inp_feat(238), I1 =>  inp_feat(505), I2 =>  inp_feat(183), I3 =>  inp_feat(365), I4 =>  inp_feat(494), I5 =>  inp_feat(30), I6 =>  inp_feat(422), I7 =>  inp_feat(362)); 
C_76_S_4_L_6_inst : LUT8 generic map(INIT => "1100111011010100110010001100100000001000100000001000100010001000010010001100000001001000110010001000100010000000100010001000100011111010100000000000101010000000001100001000000010000000100000000000101000000000000000001000000000000000000000001000000010000000") port map( O =>C_76_S_4_L_6_out, I0 =>  inp_feat(351), I1 =>  inp_feat(281), I2 =>  inp_feat(382), I3 =>  inp_feat(363), I4 =>  inp_feat(228), I5 =>  inp_feat(168), I6 =>  inp_feat(473), I7 =>  inp_feat(66)); 
C_76_S_4_L_7_inst : LUT8 generic map(INIT => "1111111111011111110110111100000011111001011110101000100000001000000100010011001100000000010100000101010110100011100000000000000000010110000010001010000000000000011100110000100000001000000000000000000000000000000000000000000001010111000000000000000000000000") port map( O =>C_76_S_4_L_7_out, I0 =>  inp_feat(478), I1 =>  inp_feat(494), I2 =>  inp_feat(388), I3 =>  inp_feat(45), I4 =>  inp_feat(426), I5 =>  inp_feat(98), I6 =>  inp_feat(381), I7 =>  inp_feat(362)); 
C_77_S_0_L_0_inst : LUT8 generic map(INIT => "1111110011101100001010101010101010000000100010101000100010001010110011001100110000000000000000000000000000000000000000000000000011101000001000000010001010101010110010100000101000000000000010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_0_L_0_out, I0 =>  inp_feat(422), I1 =>  inp_feat(381), I2 =>  inp_feat(483), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_77_S_0_L_1_inst : LUT8 generic map(INIT => "1111101011111000111100101111110011001000111000000000000000000000111000001111000000000000000000001100000010100000000000000000000010111010101100000000000000000000100000001100000000000000000000001100000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_0_L_1_out, I0 =>  inp_feat(483), I1 =>  inp_feat(78), I2 =>  inp_feat(455), I3 =>  inp_feat(422), I4 =>  inp_feat(444), I5 =>  inp_feat(338), I6 =>  inp_feat(268), I7 =>  inp_feat(505)); 
C_77_S_0_L_2_inst : LUT8 generic map(INIT => "0101110111111101111111010101000110101000111111001000000000000000111111010100011011111101110100001010000000000000100000000000000000000000100000000000000000000000100000001010000000000000000000001000000000000000100000000000000010100000000000001000000000000000") port map( O =>C_77_S_0_L_2_out, I0 =>  inp_feat(492), I1 =>  inp_feat(479), I2 =>  inp_feat(134), I3 =>  inp_feat(199), I4 =>  inp_feat(98), I5 =>  inp_feat(240), I6 =>  inp_feat(494), I7 =>  inp_feat(238)); 
C_77_S_0_L_3_inst : LUT8 generic map(INIT => "1110101010011010010000001111111110101010111001101100000000000000001000100000001010000000000000001010101000000000000000000000000011001000000000001100000000000000100010000000000010000000000000000000100000000000000000000000000000001000000000000000000000000000") port map( O =>C_77_S_0_L_3_out, I0 =>  inp_feat(134), I1 =>  inp_feat(313), I2 =>  inp_feat(240), I3 =>  inp_feat(461), I4 =>  inp_feat(432), I5 =>  inp_feat(504), I6 =>  inp_feat(281), I7 =>  inp_feat(345)); 
C_77_S_0_L_4_inst : LUT8 generic map(INIT => "1111111111111001100000000000000011111010111110110000000000000000111011001000000010000000100000001000000010000000100000001000000000000000000000000000000000000000000000001000100000000000000000000000000000000000100000001000000010000000100000001000000010000000") port map( O =>C_77_S_0_L_4_out, I0 =>  inp_feat(505), I1 =>  inp_feat(430), I2 =>  inp_feat(398), I3 =>  inp_feat(379), I4 =>  inp_feat(160), I5 =>  inp_feat(436), I6 =>  inp_feat(385), I7 =>  inp_feat(348)); 
C_77_S_0_L_5_inst : LUT8 generic map(INIT => "1110110110101101111000001010100011010000110000000000000010001000100000101110000011100010100000000000000011000000010000001000000011111101000001001111000000000000111100000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000") port map( O =>C_77_S_0_L_5_out, I0 =>  inp_feat(221), I1 =>  inp_feat(356), I2 =>  inp_feat(223), I3 =>  inp_feat(209), I4 =>  inp_feat(7), I5 =>  inp_feat(206), I6 =>  inp_feat(281), I7 =>  inp_feat(222)); 
C_77_S_0_L_6_inst : LUT8 generic map(INIT => "1111101010001000100010000000100011111010100000001010100010001000100000001000000000000000000000001100000000000000100000000000000010101010000010000000100010001000001000100000000000101010000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_0_L_6_out, I0 =>  inp_feat(160), I1 =>  inp_feat(221), I2 =>  inp_feat(430), I3 =>  inp_feat(67), I4 =>  inp_feat(338), I5 =>  inp_feat(209), I6 =>  inp_feat(237), I7 =>  inp_feat(43)); 
C_77_S_0_L_7_inst : LUT8 generic map(INIT => "1111110111111101000010000010000010000111011010111010000000101010111101011010010101010000000000001011001110101001100000101010000000000000000000000000000000000000000000000000000000001000000010001010100010100000000000000000000010100010101010000000100010000000") port map( O =>C_77_S_0_L_7_out, I0 =>  inp_feat(175), I1 =>  inp_feat(437), I2 =>  inp_feat(428), I3 =>  inp_feat(11), I4 =>  inp_feat(206), I5 =>  inp_feat(483), I6 =>  inp_feat(209), I7 =>  inp_feat(348)); 
C_77_S_1_L_0_inst : LUT8 generic map(INIT => "1111110011101100001010101010101010000000100010101000100010001010110011001100110000000000000000000000000000000000000000000000000011101000001000000010001010101010110010100000101000000000000010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_1_L_0_out, I0 =>  inp_feat(422), I1 =>  inp_feat(381), I2 =>  inp_feat(483), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_77_S_1_L_1_inst : LUT8 generic map(INIT => "1111111100101011101000001010000010101111111100110000000000000000101000000000000010100000000000000000000000000000000000000000000010100000000000000010000000000000000000000000000000000000000000001010000000000000100000000000000000000000000000000000000000000000") port map( O =>C_77_S_1_L_1_out, I0 =>  inp_feat(348), I1 =>  inp_feat(494), I2 =>  inp_feat(160), I3 =>  inp_feat(206), I4 =>  inp_feat(324), I5 =>  inp_feat(237), I6 =>  inp_feat(454), I7 =>  inp_feat(505)); 
C_77_S_1_L_2_inst : LUT8 generic map(INIT => "1111101110100010001100100000000011111111000000001111000000000000110000001100000010000000000000001100010000000000100000000000000011100010111000101100000000000000000000000000000000000000000000000000000011000000000000000000000000000000100000000000000000000000") port map( O =>C_77_S_1_L_2_out, I0 =>  inp_feat(365), I1 =>  inp_feat(235), I2 =>  inp_feat(134), I3 =>  inp_feat(313), I4 =>  inp_feat(68), I5 =>  inp_feat(72), I6 =>  inp_feat(422), I7 =>  inp_feat(240)); 
C_77_S_1_L_3_inst : LUT8 generic map(INIT => "1111101111111111111111110101011100101011100011010010101000000000110111010100010111011111010101011100110101000000000010000000000011001100000000000100000000000000000000000000000000000000000000001000110000000000100010000000000001001100000000000000000000000000") port map( O =>C_77_S_1_L_3_out, I0 =>  inp_feat(494), I1 =>  inp_feat(430), I2 =>  inp_feat(379), I3 =>  inp_feat(434), I4 =>  inp_feat(151), I5 =>  inp_feat(281), I6 =>  inp_feat(209), I7 =>  inp_feat(237)); 
C_77_S_1_L_4_inst : LUT8 generic map(INIT => "1010111110101010001010101010101000001000100000000000000010000000111111111010101010100000101010100101000000001000000000000000100010100000000000000010000010000000000000001000100000000000000000001010000010000000101000001000100000000000100010000000000010001000") port map( O =>C_77_S_1_L_4_out, I0 =>  inp_feat(455), I1 =>  inp_feat(340), I2 =>  inp_feat(7), I3 =>  inp_feat(240), I4 =>  inp_feat(351), I5 =>  inp_feat(348), I6 =>  inp_feat(494), I7 =>  inp_feat(160)); 
C_77_S_1_L_5_inst : LUT8 generic map(INIT => "1101100011111001110000000110001011001000110011110000000001100000100000101100001011000000111111110000000001001000100000001100101011101010101010100000000000000000000000000000000000000000000000001100000010000000100000001111000000000000000000000000000010010000") port map( O =>C_77_S_1_L_5_out, I0 =>  inp_feat(460), I1 =>  inp_feat(483), I2 =>  inp_feat(382), I3 =>  inp_feat(303), I4 =>  inp_feat(338), I5 =>  inp_feat(434), I6 =>  inp_feat(404), I7 =>  inp_feat(248)); 
C_77_S_1_L_6_inst : LUT8 generic map(INIT => "1111011101111110111100101111111001010010000000001111000000000000111101111101111000110000100001001101000000000000000000000000000001111111000000001111101110001000000000000000000001000000000000001101000010000000010000001000000011000000000000000000000000000000") port map( O =>C_77_S_1_L_6_out, I0 =>  inp_feat(494), I1 =>  inp_feat(88), I2 =>  inp_feat(107), I3 =>  inp_feat(358), I4 =>  inp_feat(504), I5 =>  inp_feat(381), I6 =>  inp_feat(78), I7 =>  inp_feat(390)); 
C_77_S_1_L_7_inst : LUT8 generic map(INIT => "1111101011110010111000000100000011111010111000101100000000000000010000000000000011000000000000001100000000000000010000000000000001110110011100100110110000000000111111100111001001001100000000000000110100000000100001000000000011001100000000001000100000000000") port map( O =>C_77_S_1_L_7_out, I0 =>  inp_feat(209), I1 =>  inp_feat(363), I2 =>  inp_feat(200), I3 =>  inp_feat(406), I4 =>  inp_feat(93), I5 =>  inp_feat(504), I6 =>  inp_feat(281), I7 =>  inp_feat(390)); 
C_77_S_2_L_0_inst : LUT8 generic map(INIT => "1111110011101100001010101010101010000000100010101000100010001010110011001100110000000000000000000000000000000000000000000000000011101000001000000010001010101010110010100000101000000000000010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_2_L_0_out, I0 =>  inp_feat(422), I1 =>  inp_feat(381), I2 =>  inp_feat(483), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_77_S_2_L_1_inst : LUT8 generic map(INIT => "1110110011000000100000000000000011001000100000001100000000000000111010101000000010100000101000001100101000000000000000000000000010000000000000000100000000000000110000000000000011000000000000001000100000000000000000000000000011101010000000001100000000000000") port map( O =>C_77_S_2_L_1_out, I0 =>  inp_feat(356), I1 =>  inp_feat(47), I2 =>  inp_feat(113), I3 =>  inp_feat(381), I4 =>  inp_feat(281), I5 =>  inp_feat(422), I6 =>  inp_feat(209), I7 =>  inp_feat(338)); 
C_77_S_2_L_2_inst : LUT8 generic map(INIT => "1101100011000000111000101000000011000000111000000000000000000000100000001000000011000000111100000000000010100000000000000000000011110000110100001110101011000000011000000110000000000000000000001000000011100000110000001110000001000000111000000000000010100000") port map( O =>C_77_S_2_L_2_out, I0 =>  inp_feat(434), I1 =>  inp_feat(281), I2 =>  inp_feat(160), I3 =>  inp_feat(422), I4 =>  inp_feat(209), I5 =>  inp_feat(199), I6 =>  inp_feat(338), I7 =>  inp_feat(379)); 
C_77_S_2_L_3_inst : LUT8 generic map(INIT => "0101110111011101000110001111100011011100000000000101000011110000110000000001000010000000100000001100000000000000110100001111000010011000100010001011100010001000110011000000000001010000010100001000000010000000000000001000000001000000000000001100000001000000") port map( O =>C_77_S_2_L_3_out, I0 =>  inp_feat(399), I1 =>  inp_feat(256), I2 =>  inp_feat(345), I3 =>  inp_feat(166), I4 =>  inp_feat(11), I5 =>  inp_feat(358), I6 =>  inp_feat(328), I7 =>  inp_feat(102)); 
C_77_S_2_L_4_inst : LUT8 generic map(INIT => "1110100011001100101010001100100010001000100000001000100011001100111000001100110011100000000000001100100011001100111010001100100000000000000000001000000000000000000000000000000000000000000000001011000000000000111000000000000000000000000000000010000000000000") port map( O =>C_77_S_2_L_4_out, I0 =>  inp_feat(167), I1 =>  inp_feat(160), I2 =>  inp_feat(355), I3 =>  inp_feat(199), I4 =>  inp_feat(379), I5 =>  inp_feat(352), I6 =>  inp_feat(240), I7 =>  inp_feat(348)); 
C_77_S_2_L_5_inst : LUT8 generic map(INIT => "1111110011001110111110000000000011011100100011001000000000000000111010001010101011000000000000001100000000000000110000000000000000001010000010000000000000000000000000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000") port map( O =>C_77_S_2_L_5_out, I0 =>  inp_feat(199), I1 =>  inp_feat(194), I2 =>  inp_feat(388), I3 =>  inp_feat(238), I4 =>  inp_feat(134), I5 =>  inp_feat(479), I6 =>  inp_feat(334), I7 =>  inp_feat(79)); 
C_77_S_2_L_6_inst : LUT8 generic map(INIT => "1111111111000100111110001110000011111111110000001111110000100000110000000000000000000000000000001000100000000000000010000000000011011010000000001111100000000000111111010000000001110000000000001100000000000000100000000000000000000000000000000000000000000000") port map( O =>C_77_S_2_L_6_out, I0 =>  inp_feat(460), I1 =>  inp_feat(479), I2 =>  inp_feat(338), I3 =>  inp_feat(455), I4 =>  inp_feat(190), I5 =>  inp_feat(265), I6 =>  inp_feat(206), I7 =>  inp_feat(483)); 
C_77_S_2_L_7_inst : LUT8 generic map(INIT => "1111110010100000111111101000100011000000100000001100000010001000110000000000000011100000000000001110000011000000111000001100000010001100000000001111110100000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_2_L_7_out, I0 =>  inp_feat(298), I1 =>  inp_feat(281), I2 =>  inp_feat(245), I3 =>  inp_feat(25), I4 =>  inp_feat(494), I5 =>  inp_feat(125), I6 =>  inp_feat(381), I7 =>  inp_feat(461)); 
C_77_S_3_L_0_inst : LUT8 generic map(INIT => "1111110011101100001010101010101010000000100010101000100010001010110011001100110000000000000000000000000000000000000000000000000011101000001000000010001010101010110010100000101000000000000010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_3_L_0_out, I0 =>  inp_feat(422), I1 =>  inp_feat(381), I2 =>  inp_feat(483), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_77_S_3_L_1_inst : LUT8 generic map(INIT => "1110110011000000100000000000000011001000100000001100000000000000111010101000000010100000101000001100101000000000000000000000000010000000000000000100000000000000110000000000000011000000000000001000100000000000000000000000000011101010000000001100000000000000") port map( O =>C_77_S_3_L_1_out, I0 =>  inp_feat(356), I1 =>  inp_feat(47), I2 =>  inp_feat(113), I3 =>  inp_feat(381), I4 =>  inp_feat(281), I5 =>  inp_feat(422), I6 =>  inp_feat(209), I7 =>  inp_feat(338)); 
C_77_S_3_L_2_inst : LUT8 generic map(INIT => "1111111011100000000000000000000011000100000000001100000000000000110011000000000000001000000000001100010000000000000010000000000011101110111000001100100000000000110001000000000000000000000000001100110000000000000010000000000001001100000000000000100000000000") port map( O =>C_77_S_3_L_2_out, I0 =>  inp_feat(171), I1 =>  inp_feat(206), I2 =>  inp_feat(324), I3 =>  inp_feat(237), I4 =>  inp_feat(454), I5 =>  inp_feat(505), I6 =>  inp_feat(199), I7 =>  inp_feat(379)); 
C_77_S_3_L_3_inst : LUT8 generic map(INIT => "0001100011001000010110000010000011010010100010000001000000010000110101011110000011111001000000000101010100000000010101010000000011011001100010101111001000110010110010101010101000010000001000101101010110101010110111010000000000001000101010100000000000000000") port map( O =>C_77_S_3_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(461), I2 =>  inp_feat(430), I3 =>  inp_feat(50), I4 =>  inp_feat(221), I5 =>  inp_feat(3), I6 =>  inp_feat(494), I7 =>  inp_feat(88)); 
C_77_S_3_L_4_inst : LUT8 generic map(INIT => "1111110000001000100000000000000011101000101010001110100010101000110111010000000010001000000000001010000000000000100000000000000011000000000000001000000000000000100000000000000010000000100000000100000000000000000000000000000010100000000000001000000000000000") port map( O =>C_77_S_3_L_4_out, I0 =>  inp_feat(298), I1 =>  inp_feat(79), I2 =>  inp_feat(483), I3 =>  inp_feat(348), I4 =>  inp_feat(238), I5 =>  inp_feat(209), I6 =>  inp_feat(406), I7 =>  inp_feat(194)); 
C_77_S_3_L_5_inst : LUT8 generic map(INIT => "1101100010001000110010000000000011111000110100001100100000000000111110000000000011001000000000001111000001110000110011000000000010001000000000001000000000000000000010000000000010001000000000000000110000000000100010000000000000000000000000000000000000000000") port map( O =>C_77_S_3_L_5_out, I0 =>  inp_feat(72), I1 =>  inp_feat(455), I2 =>  inp_feat(135), I3 =>  inp_feat(237), I4 =>  inp_feat(343), I5 =>  inp_feat(359), I6 =>  inp_feat(298), I7 =>  inp_feat(248)); 
C_77_S_3_L_6_inst : LUT8 generic map(INIT => "1101110011001000111111001000100001000000100010001111100010101010110011001000000011000000000000000000000000000000110000000000000011001100100000001100000000000000100000001000000011000000000000000100000010000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_3_L_6_out, I0 =>  inp_feat(135), I1 =>  inp_feat(348), I2 =>  inp_feat(194), I3 =>  inp_feat(171), I4 =>  inp_feat(209), I5 =>  inp_feat(238), I6 =>  inp_feat(298), I7 =>  inp_feat(356)); 
C_77_S_3_L_7_inst : LUT8 generic map(INIT => "1101110011011100100010001000000010001100110010001100000011000000100110001111110010001000000000000000100000000000100000001000000010100100010010001000000011000000110010001100000000000000110000001111110011001100110000000100000000000000000000001000000000000000") port map( O =>C_77_S_3_L_7_out, I0 =>  inp_feat(80), I1 =>  inp_feat(348), I2 =>  inp_feat(338), I3 =>  inp_feat(468), I4 =>  inp_feat(221), I5 =>  inp_feat(318), I6 =>  inp_feat(135), I7 =>  inp_feat(483)); 
C_77_S_4_L_0_inst : LUT8 generic map(INIT => "1111110011101100001010101010101010000000100010101000100010001010110011001100110000000000000000000000000000000000000000000000000011101000001000000010001010101010110010100000101000000000000010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_4_L_0_out, I0 =>  inp_feat(422), I1 =>  inp_feat(381), I2 =>  inp_feat(483), I3 =>  inp_feat(494), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_77_S_4_L_1_inst : LUT8 generic map(INIT => "1110110011001000110000001000000010000000110000000000000000000000111010101100101010000000000000001010000000000000101000000000000010000000110000000000000000000000010000001100000000000000000000001000100011101010000000000000000000000000110000000000000000000000") port map( O =>C_77_S_4_L_1_out, I0 =>  inp_feat(356), I1 =>  inp_feat(47), I2 =>  inp_feat(113), I3 =>  inp_feat(422), I4 =>  inp_feat(381), I5 =>  inp_feat(281), I6 =>  inp_feat(209), I7 =>  inp_feat(338)); 
C_77_S_4_L_2_inst : LUT8 generic map(INIT => "1111111011100000000000000000000011000100000000001100000000000000110011000000000000001000000000001100010000000000000010000000000011101110111000001100100000000000110001000000000000000000000000001100110000000000000010000000000001001100000000000000100000000000") port map( O =>C_77_S_4_L_2_out, I0 =>  inp_feat(171), I1 =>  inp_feat(206), I2 =>  inp_feat(324), I3 =>  inp_feat(237), I4 =>  inp_feat(454), I5 =>  inp_feat(505), I6 =>  inp_feat(199), I7 =>  inp_feat(379)); 
C_77_S_4_L_3_inst : LUT8 generic map(INIT => "0001100011001000010110000010000011010010100010000001000000010000110101011110000011111001000000000101010100000000010101010000000011011001100010101111001000110010110010101010101000010000001000101101010110101010110111010000000000001000101010100000000000000000") port map( O =>C_77_S_4_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(461), I2 =>  inp_feat(430), I3 =>  inp_feat(50), I4 =>  inp_feat(221), I5 =>  inp_feat(3), I6 =>  inp_feat(494), I7 =>  inp_feat(88)); 
C_77_S_4_L_4_inst : LUT8 generic map(INIT => "1111110000001000100000000000000011101000101010001110100010101000110111010000000010001000000000001010000000000000100000000000000011000000000000001000000000000000100000000000000010000000100000000100000000000000000000000000000010100000000000001000000000000000") port map( O =>C_77_S_4_L_4_out, I0 =>  inp_feat(298), I1 =>  inp_feat(79), I2 =>  inp_feat(483), I3 =>  inp_feat(348), I4 =>  inp_feat(238), I5 =>  inp_feat(209), I6 =>  inp_feat(406), I7 =>  inp_feat(194)); 
C_77_S_4_L_5_inst : LUT8 generic map(INIT => "1101100010001000110010000000000011111000110100001100100000000000111110000000000011001000000000001111000001110000110011000000000010001000000000001000000000000000000010000000000010001000000000000000110000000000100010000000000000000000000000000000000000000000") port map( O =>C_77_S_4_L_5_out, I0 =>  inp_feat(72), I1 =>  inp_feat(455), I2 =>  inp_feat(135), I3 =>  inp_feat(237), I4 =>  inp_feat(343), I5 =>  inp_feat(359), I6 =>  inp_feat(298), I7 =>  inp_feat(248)); 
C_77_S_4_L_6_inst : LUT8 generic map(INIT => "1101110011001000111111001000100001000000100010001111100010101010110011001000000011000000000000000000000000000000110000000000000011001100100000001100000000000000100000001000000011000000000000000100000010000000000000000000000000000000000000000000000000000000") port map( O =>C_77_S_4_L_6_out, I0 =>  inp_feat(135), I1 =>  inp_feat(348), I2 =>  inp_feat(194), I3 =>  inp_feat(171), I4 =>  inp_feat(209), I5 =>  inp_feat(238), I6 =>  inp_feat(298), I7 =>  inp_feat(356)); 
C_77_S_4_L_7_inst : LUT8 generic map(INIT => "1101110011011100100010001000000010001100110010001100000011000000100110001111110010001000000000000000100000000000100000001000000010100100010010001000000011000000110010001100000000000000110000001111110011001100110000000100000000000000000000001000000000000000") port map( O =>C_77_S_4_L_7_out, I0 =>  inp_feat(80), I1 =>  inp_feat(348), I2 =>  inp_feat(338), I3 =>  inp_feat(468), I4 =>  inp_feat(221), I5 =>  inp_feat(318), I6 =>  inp_feat(135), I7 =>  inp_feat(483)); 
C_78_S_0_L_0_inst : LUT8 generic map(INIT => "1110111110100000111001001110110011001111000100001100111101100010111000001010000010100000101000001000000000000000000000000000000011001101100000001010010100000000110011100000000010001110000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_78_S_0_L_0_out, I0 =>  inp_feat(259), I1 =>  inp_feat(342), I2 =>  inp_feat(502), I3 =>  inp_feat(256), I4 =>  inp_feat(469), I5 =>  inp_feat(330), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_78_S_0_L_1_inst : LUT8 generic map(INIT => "0001011100010111111111110001111100100000111000000000000010000000000100000000001011100011011000100000000010000000101000001000000011010101110000001000000010000000010000001100000000000000100000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_78_S_0_L_1_out, I0 =>  inp_feat(98), I1 =>  inp_feat(184), I2 =>  inp_feat(126), I3 =>  inp_feat(77), I4 =>  inp_feat(178), I5 =>  inp_feat(461), I6 =>  inp_feat(202), I7 =>  inp_feat(242)); 
C_78_S_0_L_2_inst : LUT8 generic map(INIT => "0000000000001000001011000000000000000000000000000000000000000000110010100010101010001011010010111110101010001010110000000000000011001000000000001100000000000000100000001000000010000000000000001000100000000000000000000000000010001000100000001000000010000000") port map( O =>C_78_S_0_L_2_out, I0 =>  inp_feat(74), I1 =>  inp_feat(238), I2 =>  inp_feat(93), I3 =>  inp_feat(21), I4 =>  inp_feat(149), I5 =>  inp_feat(116), I6 =>  inp_feat(494), I7 =>  inp_feat(492)); 
C_78_S_0_L_3_inst : LUT8 generic map(INIT => "0011110010100000110111111000100000000000000000001000100010000000001111101100110011011111101010100000000010000000100010101000100000111000000000001111101000111011000000000000000000111010001100110010000000000010101000101000101000000000000000000000000010100010") port map( O =>C_78_S_0_L_3_out, I0 =>  inp_feat(149), I1 =>  inp_feat(30), I2 =>  inp_feat(420), I3 =>  inp_feat(164), I4 =>  inp_feat(494), I5 =>  inp_feat(339), I6 =>  inp_feat(331), I7 =>  inp_feat(114)); 
C_78_S_0_L_4_inst : LUT8 generic map(INIT => "1111110000001111101011100000111100011000001101001110100100010100111011001000000010001100000000001000100000000000100011001000000000001000000010000000111000000000000000000000000000000110000000001111111110100000101000001010000001000100100000000000100010100000") port map( O =>C_78_S_0_L_4_out, I0 =>  inp_feat(259), I1 =>  inp_feat(383), I2 =>  inp_feat(365), I3 =>  inp_feat(449), I4 =>  inp_feat(475), I5 =>  inp_feat(362), I6 =>  inp_feat(102), I7 =>  inp_feat(370)); 
C_78_S_0_L_5_inst : LUT8 generic map(INIT => "0101111011111001111110010100010000111000111111000011000101010100111100000101010011111010110111011111000001000000100010011101110100101000001110001100000011111111000000000010000001110001011100011111000011111000111010011111111100001000010100101001100011111111") port map( O =>C_78_S_0_L_5_out, I0 =>  inp_feat(468), I1 =>  inp_feat(340), I2 =>  inp_feat(440), I3 =>  inp_feat(98), I4 =>  inp_feat(276), I5 =>  inp_feat(190), I6 =>  inp_feat(219), I7 =>  inp_feat(110)); 
C_78_S_0_L_6_inst : LUT8 generic map(INIT => "0101001010100010011101001111010010101000101010101111110111111110011100001010000000110100010001000000000000000000000000000000010010100000100000000010000010000000000010001000000010110010111100101010000000000000000000000000000000000000000000000000000000000000") port map( O =>C_78_S_0_L_6_out, I0 =>  inp_feat(30), I1 =>  inp_feat(31), I2 =>  inp_feat(261), I3 =>  inp_feat(420), I4 =>  inp_feat(58), I5 =>  inp_feat(228), I6 =>  inp_feat(80), I7 =>  inp_feat(271)); 
C_78_S_0_L_7_inst : LUT8 generic map(INIT => "1110110010000000111010000010000011101010011000100010000000100000111011011000000011110111110000010000010101010101000100011111010110000000000000001000000000100000101010000000000000000000001000001100110000000000101010000000000010001000000000000000100000000000") port map( O =>C_78_S_0_L_7_out, I0 =>  inp_feat(344), I1 =>  inp_feat(491), I2 =>  inp_feat(206), I3 =>  inp_feat(250), I4 =>  inp_feat(65), I5 =>  inp_feat(95), I6 =>  inp_feat(316), I7 =>  inp_feat(114)); 
C_78_S_1_L_0_inst : LUT8 generic map(INIT => "1111101010111010111110111111100010110000000000000111000000000000111110001111000011111000110100001111000011010000010100000000000000100000101000100010000011100000000000000000000000000000000000000100000000000000010000000000000000100000000000000000000000000000") port map( O =>C_78_S_1_L_0_out, I0 =>  inp_feat(323), I1 =>  inp_feat(340), I2 =>  inp_feat(193), I3 =>  inp_feat(289), I4 =>  inp_feat(290), I5 =>  inp_feat(190), I6 =>  inp_feat(125), I7 =>  inp_feat(80)); 
C_78_S_1_L_1_inst : LUT8 generic map(INIT => "1100101011011000000010001000100010101000100010101000100000001000111011101100110011011101000011011110110011011101010011001100110110000010010010100000000000100100000010000000101100000000100011111000111000000101100110000000010110101100110011011100110000001101") port map( O =>C_78_S_1_L_1_out, I0 =>  inp_feat(409), I1 =>  inp_feat(281), I2 =>  inp_feat(7), I3 =>  inp_feat(401), I4 =>  inp_feat(362), I5 =>  inp_feat(93), I6 =>  inp_feat(494), I7 =>  inp_feat(80)); 
C_78_S_1_L_2_inst : LUT8 generic map(INIT => "1110000100101100100000001010000010101010111010001010100011101100000000000000000000000000001000000010000000100000000000000010000011111000100000001000100010111000111010001000100010001000100010001010000000000000100010000000000000000000000000001000100010001000") port map( O =>C_78_S_1_L_2_out, I0 =>  inp_feat(114), I1 =>  inp_feat(426), I2 =>  inp_feat(362), I3 =>  inp_feat(492), I4 =>  inp_feat(61), I5 =>  inp_feat(170), I6 =>  inp_feat(502), I7 =>  inp_feat(89)); 
C_78_S_1_L_3_inst : LUT8 generic map(INIT => "1111110111110110111111011111010011100111001100001111010100000000101011101110000011000000001100000010000000100000011001000000000001000100000001001100000000000000010001000000000000000000000000001110111000000000000000000000000000000100000000000000000000000000") port map( O =>C_78_S_1_L_3_out, I0 =>  inp_feat(340), I1 =>  inp_feat(437), I2 =>  inp_feat(406), I3 =>  inp_feat(374), I4 =>  inp_feat(249), I5 =>  inp_feat(356), I6 =>  inp_feat(396), I7 =>  inp_feat(190)); 
C_78_S_1_L_4_inst : LUT8 generic map(INIT => "1011101011101101000000001000100010111110111111100000000010000000101010110000000000100000000000001000111110100000101100001111000010100011000001000000100000000000000110100001000100000000000000000010001000000000000000000000000000001111000000000000101100010000") port map( O =>C_78_S_1_L_4_out, I0 =>  inp_feat(105), I1 =>  inp_feat(247), I2 =>  inp_feat(65), I3 =>  inp_feat(494), I4 =>  inp_feat(319), I5 =>  inp_feat(420), I6 =>  inp_feat(358), I7 =>  inp_feat(181)); 
C_78_S_1_L_5_inst : LUT8 generic map(INIT => "0011001010110101111111101010010010001100000011001000100010000101111111001111111111001111111011110000000001110010100000110100111100111100001100010100000101100000000010001100000000000101010001111000000011100011000000001111011100001000111101111000110111111111") port map( O =>C_78_S_1_L_5_out, I0 =>  inp_feat(120), I1 =>  inp_feat(477), I2 =>  inp_feat(504), I3 =>  inp_feat(388), I4 =>  inp_feat(259), I5 =>  inp_feat(77), I6 =>  inp_feat(330), I7 =>  inp_feat(238)); 
C_78_S_1_L_6_inst : LUT8 generic map(INIT => "1101010110001101100101011101110101111111110111010101110100000101000100001000100000000000100010000101010111010101000101010000100101111101110110010001010100010000111111110101110101010101000101010001000000000000000000000000000000000001010101010001000100010101") port map( O =>C_78_S_1_L_6_out, I0 =>  inp_feat(170), I1 =>  inp_feat(475), I2 =>  inp_feat(431), I3 =>  inp_feat(45), I4 =>  inp_feat(66), I5 =>  inp_feat(358), I6 =>  inp_feat(237), I7 =>  inp_feat(473)); 
C_78_S_1_L_7_inst : LUT8 generic map(INIT => "0111111000000000000000000010000001110100011111001100000000001100010011010000101010001000000000101100110011111111110000000101110111001111100011011011111101011111000011001001111101000000011111110100110000001100010010000001011100001110000011110000110111111101") port map( O =>C_78_S_1_L_7_out, I0 =>  inp_feat(492), I1 =>  inp_feat(459), I2 =>  inp_feat(219), I3 =>  inp_feat(486), I4 =>  inp_feat(137), I5 =>  inp_feat(170), I6 =>  inp_feat(268), I7 =>  inp_feat(311)); 
C_78_S_2_L_0_inst : LUT8 generic map(INIT => "1101110111110000000010101010101010011100111111111000110000001000100011101000000000001111000000001100110001001100000010000000000011000100110001000000001000101010110011001100110000001000100010000000000000000100000000000000000000000100110001000000000000000000") port map( O =>C_78_S_2_L_0_out, I0 =>  inp_feat(468), I1 =>  inp_feat(357), I2 =>  inp_feat(102), I3 =>  inp_feat(170), I4 =>  inp_feat(508), I5 =>  inp_feat(312), I6 =>  inp_feat(502), I7 =>  inp_feat(268)); 
C_78_S_2_L_1_inst : LUT8 generic map(INIT => "0100110011001000001010100000000011100000110000000010000000000000011010111100011110101010100000000000000000000010000000000000000011111111111101010101010100000000111111110001000000010000000000001011101111111111111100010011101100010011011101110100000000000000") port map( O =>C_78_S_2_L_1_out, I0 =>  inp_feat(492), I1 =>  inp_feat(102), I2 =>  inp_feat(85), I3 =>  inp_feat(57), I4 =>  inp_feat(508), I5 =>  inp_feat(502), I6 =>  inp_feat(268), I7 =>  inp_feat(312)); 
C_78_S_2_L_2_inst : LUT8 generic map(INIT => "1100110111100000010000001100100011001100110000000000100011000000000010000100000000000000000000001100100000000000110000000000000001001100000000000000000001000000011101100100000000000000110000000000000000000000000000000000000011000000000000000000000000000000") port map( O =>C_78_S_2_L_2_out, I0 =>  inp_feat(290), I1 =>  inp_feat(348), I2 =>  inp_feat(270), I3 =>  inp_feat(241), I4 =>  inp_feat(451), I5 =>  inp_feat(161), I6 =>  inp_feat(190), I7 =>  inp_feat(80)); 
C_78_S_2_L_3_inst : LUT8 generic map(INIT => "1011001101110111011111110000010111100000101000000010000000000000101111111001111101001111010011111110001010101010000000100000101011010000000000011101010000010000111000000000000010010010000001111111101100011111110001010001000010100101000010110000010101000001") port map( O =>C_78_S_2_L_3_out, I0 =>  inp_feat(388), I1 =>  inp_feat(120), I2 =>  inp_feat(502), I3 =>  inp_feat(149), I4 =>  inp_feat(21), I5 =>  inp_feat(161), I6 =>  inp_feat(270), I7 =>  inp_feat(77)); 
C_78_S_2_L_4_inst : LUT8 generic map(INIT => "0001101101111111001011001011001110000010101000101110000010000010100010001110101011000000111000101100000011000000110000001110000011101000110010100010000000000000111000001100000000100000000000001000000011000000000000000000000011000000110000000000000000000000") port map( O =>C_78_S_2_L_4_out, I0 =>  inp_feat(362), I1 =>  inp_feat(312), I2 =>  inp_feat(493), I3 =>  inp_feat(420), I4 =>  inp_feat(396), I5 =>  inp_feat(470), I6 =>  inp_feat(152), I7 =>  inp_feat(394)); 
C_78_S_2_L_5_inst : LUT8 generic map(INIT => "1111001001001100010011111000110000010001000101000000000000000100111111101000000001001101100000000000000000000000000000000000000011111100110011100000010000000100111000000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000") port map( O =>C_78_S_2_L_5_out, I0 =>  inp_feat(102), I1 =>  inp_feat(398), I2 =>  inp_feat(374), I3 =>  inp_feat(401), I4 =>  inp_feat(76), I5 =>  inp_feat(281), I6 =>  inp_feat(24), I7 =>  inp_feat(431)); 
C_78_S_2_L_6_inst : LUT8 generic map(INIT => "1011111100101111000101000010111111011101110111111111110111111111101111001111110001010000010000001100010000000101000000000001000011001001100000000000000010000000000000001101010000010000111100011000100010000001100100000001000100000000000001010001000000000001") port map( O =>C_78_S_2_L_6_out, I0 =>  inp_feat(232), I1 =>  inp_feat(303), I2 =>  inp_feat(346), I3 =>  inp_feat(277), I4 =>  inp_feat(238), I5 =>  inp_feat(330), I6 =>  inp_feat(131), I7 =>  inp_feat(342)); 
C_78_S_2_L_7_inst : LUT8 generic map(INIT => "0111011101110001000000011111110010000110100000001100111100000000010001111101101000001101110101110000000001000100000001110000001101101110110011000101110101011101000011000000000011000111000001110000000011001100010101110110001000000000010001000000011101011111") port map( O =>C_78_S_2_L_7_out, I0 =>  inp_feat(309), I1 =>  inp_feat(412), I2 =>  inp_feat(388), I3 =>  inp_feat(232), I4 =>  inp_feat(307), I5 =>  inp_feat(271), I6 =>  inp_feat(100), I7 =>  inp_feat(93)); 
C_78_S_3_L_0_inst : LUT8 generic map(INIT => "1011110011110000011100010111001111100000110000000000000000000000111011001010000010100100101000001100110000000000000000000000000000000000110000000000000000110010000000000000000000000000010000001000100000000000100001000000000000000000000000000000010000000000") port map( O =>C_78_S_3_L_0_out, I0 =>  inp_feat(102), I1 =>  inp_feat(276), I2 =>  inp_feat(502), I3 =>  inp_feat(312), I4 =>  inp_feat(68), I5 =>  inp_feat(342), I6 =>  inp_feat(250), I7 =>  inp_feat(507)); 
C_78_S_3_L_1_inst : LUT8 generic map(INIT => "0010000000000000101000000000000011101100110001010111101000110000101000100100111000000000000000001010001011001110000000000000000011101111110000001011110010000000101011100000000000000010000000000100101111001111010000001100000000001010000011110000000000000000") port map( O =>C_78_S_3_L_1_out, I0 =>  inp_feat(362), I1 =>  inp_feat(505), I2 =>  inp_feat(43), I3 =>  inp_feat(413), I4 =>  inp_feat(74), I5 =>  inp_feat(396), I6 =>  inp_feat(414), I7 =>  inp_feat(494)); 
C_78_S_3_L_2_inst : LUT8 generic map(INIT => "1110011101101000010111000100110101010001000000000000010000000000111011111110000001100101011100001101111100000000100000010000000011001110110011000000000101000100000000000000000000000000000000001101010111000100010101010000000011010101000000000101000100000000") port map( O =>C_78_S_3_L_2_out, I0 =>  inp_feat(95), I1 =>  inp_feat(306), I2 =>  inp_feat(340), I3 =>  inp_feat(259), I4 =>  inp_feat(440), I5 =>  inp_feat(268), I6 =>  inp_feat(471), I7 =>  inp_feat(24)); 
C_78_S_3_L_3_inst : LUT8 generic map(INIT => "0101111100001100101010001000100001101111000001000000000000001000111101110000000010100000000000000100011100000000000000000000000011000000100000001000100010101000101000001010101000101000101010101000100000000000101010101010100010100011100000001010101010101010") port map( O =>C_78_S_3_L_3_out, I0 =>  inp_feat(312), I1 =>  inp_feat(6), I2 =>  inp_feat(309), I3 =>  inp_feat(390), I4 =>  inp_feat(363), I5 =>  inp_feat(100), I6 =>  inp_feat(378), I7 =>  inp_feat(70)); 
C_78_S_3_L_4_inst : LUT8 generic map(INIT => "1111110011101110101000001110111010111000110011001010000000000000000000001100110100000010111010010000000000000000001000000000000011100010110011001110001011001100000010001100100000100000110011001000101000000000101010101100110000001000010000001010110011001100") port map( O =>C_78_S_3_L_4_out, I0 =>  inp_feat(383), I1 =>  inp_feat(413), I2 =>  inp_feat(80), I3 =>  inp_feat(404), I4 =>  inp_feat(379), I5 =>  inp_feat(461), I6 =>  inp_feat(281), I7 =>  inp_feat(296)); 
C_78_S_3_L_5_inst : LUT8 generic map(INIT => "0111111011010010110101101100001011110111011001101101011110001111011010101010001001000010010000101110001000100010000000000010001011011111010100100111111101001000000101110000000001011100011101011110001000000010010000100100000000100010001000100000000000100010") port map( O =>C_78_S_3_L_5_out, I0 =>  inp_feat(492), I1 =>  inp_feat(508), I2 =>  inp_feat(385), I3 =>  inp_feat(100), I4 =>  inp_feat(6), I5 =>  inp_feat(486), I6 =>  inp_feat(475), I7 =>  inp_feat(378)); 
C_78_S_3_L_6_inst : LUT8 generic map(INIT => "0011010110110001111100001000000111110011001000101111000100100000100110011000101000110100111101110011010111111111001100000011001111110010001100101111000000000000000100000010000000110000000000000001001100000001111100011101010111110010010111110111001000010000") port map( O =>C_78_S_3_L_6_out, I0 =>  inp_feat(98), I1 =>  inp_feat(388), I2 =>  inp_feat(237), I3 =>  inp_feat(149), I4 =>  inp_feat(263), I5 =>  inp_feat(477), I6 =>  inp_feat(344), I7 =>  inp_feat(357)); 
C_78_S_3_L_7_inst : LUT8 generic map(INIT => "1100001111001101101010010000010010101111110000001111110110101110111010101100111110001100110111111000110010101111111011111110111100000100000011001100100010001000000000001000100001110000001010000000100000000110000000000010000000001100101011100000000010101111") port map( O =>C_78_S_3_L_7_out, I0 =>  inp_feat(238), I1 =>  inp_feat(263), I2 =>  inp_feat(388), I3 =>  inp_feat(129), I4 =>  inp_feat(27), I5 =>  inp_feat(259), I6 =>  inp_feat(330), I7 =>  inp_feat(357)); 
C_78_S_4_L_0_inst : LUT8 generic map(INIT => "1010001010100101111110001000000111100100001000001100110000100000111110001110000010000000111010000010000001100000000000001110000011011100000010001111110001111101111111001100110101101100001000001110100011110100101000001111110111101000111001100010000011111111") port map( O =>C_78_S_4_L_0_out, I0 =>  inp_feat(468), I1 =>  inp_feat(351), I2 =>  inp_feat(362), I3 =>  inp_feat(507), I4 =>  inp_feat(493), I5 =>  inp_feat(100), I6 =>  inp_feat(93), I7 =>  inp_feat(3)); 
C_78_S_4_L_1_inst : LUT8 generic map(INIT => "1100010010011101110111001101110011000001010100001101110010000100111100011101010111111101110111010101110100001101111111111101111111100000111100001000100000000000000000000000000000000000000000001111100011110011110110010101011100000100011011110101110101011111") port map( O =>C_78_S_4_L_1_out, I0 =>  inp_feat(492), I1 =>  inp_feat(502), I2 =>  inp_feat(85), I3 =>  inp_feat(459), I4 =>  inp_feat(219), I5 =>  inp_feat(268), I6 =>  inp_feat(471), I7 =>  inp_feat(24)); 
C_78_S_4_L_2_inst : LUT8 generic map(INIT => "0100111001111100110011111101110011111111000001001011111111011100000011100001000001010000010001000100000000010001100000000001010010001101100011001000100010001100100010000000000010000000000011000000000000000000000010000000100000000000000000000000000000000000") port map( O =>C_78_S_4_L_2_out, I0 =>  inp_feat(504), I1 =>  inp_feat(413), I2 =>  inp_feat(328), I3 =>  inp_feat(216), I4 =>  inp_feat(494), I5 =>  inp_feat(460), I6 =>  inp_feat(238), I7 =>  inp_feat(262)); 
C_78_S_4_L_3_inst : LUT8 generic map(INIT => "1111011111111111111011111111111111111000111110101000000101001000111010101010101011100010000010100111000010111010000000001000101000000111010101000000000001010010000100000000000000000000000000000010000010101010000000001010101000000000100010100000000000000000") port map( O =>C_78_S_4_L_3_out, I0 =>  inp_feat(396), I1 =>  inp_feat(87), I2 =>  inp_feat(135), I3 =>  inp_feat(493), I4 =>  inp_feat(383), I5 =>  inp_feat(461), I6 =>  inp_feat(296), I7 =>  inp_feat(281)); 
C_78_S_4_L_4_inst : LUT8 generic map(INIT => "0100101011001000111010101100110000000010110000001110010010001000100010001000100000100010000000000000000000000000000000100000000011001100010101001111111111101111000011000000000000001010000000001001010100000100011101110111111000000000000000000000001000000000") port map( O =>C_78_S_4_L_4_out, I0 =>  inp_feat(100), I1 =>  inp_feat(237), I2 =>  inp_feat(385), I3 =>  inp_feat(378), I4 =>  inp_feat(98), I5 =>  inp_feat(95), I6 =>  inp_feat(47), I7 =>  inp_feat(70)); 
C_78_S_4_L_5_inst : LUT8 generic map(INIT => "1110011010101000110110011011111110100000100000000010000010110111101000000000000010100010000000001010001000000000001000000000000010001010100010001010001010101000001000000000000000100000000000000000001000000000001000100000000000000000000000000000000000000000") port map( O =>C_78_S_4_L_5_out, I0 =>  inp_feat(441), I1 =>  inp_feat(350), I2 =>  inp_feat(459), I3 =>  inp_feat(24), I4 =>  inp_feat(93), I5 =>  inp_feat(137), I6 =>  inp_feat(281), I7 =>  inp_feat(383)); 
C_78_S_4_L_6_inst : LUT8 generic map(INIT => "0110011110001111000001110000010111011111000110111000011100010100111101110011001101101011001101111011011100110011001110110011001111111111001101110011111100000001111111110100000100001111000000001111111100110011011111110001001100110011000100110011001100000011") port map( O =>C_78_S_4_L_6_out, I0 =>  inp_feat(120), I1 =>  inp_feat(277), I2 =>  inp_feat(98), I3 =>  inp_feat(462), I4 =>  inp_feat(357), I5 =>  inp_feat(263), I6 =>  inp_feat(393), I7 =>  inp_feat(477)); 
C_78_S_4_L_7_inst : LUT8 generic map(INIT => "1100100011111111110010001101010010100000100000010000000010000001110100001110110111001100110001010000000010101000000001001010010110100000100101010000000000000000101001110010001100000000000001010110100111101101000000000000100001100000011011010101010001010100") port map( O =>C_78_S_4_L_7_out, I0 =>  inp_feat(105), I1 =>  inp_feat(351), I2 =>  inp_feat(295), I3 =>  inp_feat(494), I4 =>  inp_feat(21), I5 =>  inp_feat(280), I6 =>  inp_feat(177), I7 =>  inp_feat(30)); 
C_79_S_0_L_0_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000001010100000000001100110000000000000011000000000001000000000000000100111000000000") port map( O =>C_79_S_0_L_0_out, I0 =>  inp_feat(23), I1 =>  inp_feat(95), I2 =>  inp_feat(68), I3 =>  inp_feat(141), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_79_S_0_L_1_inst : LUT8 generic map(INIT => "0010000000010000000000000000000000000001000000100000100100001000000000000001000000000000000000000000100000001011000000000000000100000000000000000000000001000100000000001010111100000000000011010000000000000000000000000000000000000010000010110000001000000010") port map( O =>C_79_S_0_L_1_out, I0 =>  inp_feat(372), I1 =>  inp_feat(348), I2 =>  inp_feat(160), I3 =>  inp_feat(338), I4 =>  inp_feat(47), I5 =>  inp_feat(194), I6 =>  inp_feat(451), I7 =>  inp_feat(505)); 
C_79_S_0_L_2_inst : LUT8 generic map(INIT => "1011101000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_0_L_2_out, I0 =>  inp_feat(27), I1 =>  inp_feat(206), I2 =>  inp_feat(467), I3 =>  inp_feat(88), I4 =>  inp_feat(170), I5 =>  inp_feat(326), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_79_S_0_L_3_inst : LUT8 generic map(INIT => "0000000000100000001100000011000000000000001000001000000000110000000000000000000000000000000000000000000000000000010000000000000000000000100000000001000010110000000000000000000000000000001000000000000000000000000000001010000000000000000000000000000000000000") port map( O =>C_79_S_0_L_3_out, I0 =>  inp_feat(468), I1 =>  inp_feat(190), I2 =>  inp_feat(399), I3 =>  inp_feat(245), I4 =>  inp_feat(281), I5 =>  inp_feat(215), I6 =>  inp_feat(95), I7 =>  inp_feat(377)); 
C_79_S_0_L_4_inst : LUT8 generic map(INIT => "1000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_0_L_4_out, I0 =>  inp_feat(170), I1 =>  inp_feat(504), I2 =>  inp_feat(47), I3 =>  inp_feat(228), I4 =>  inp_feat(88), I5 =>  inp_feat(92), I6 =>  inp_feat(209), I7 =>  inp_feat(72)); 
C_79_S_0_L_5_inst : LUT8 generic map(INIT => "0000000001000000011100100000000001110010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_0_L_5_out, I0 =>  inp_feat(145), I1 =>  inp_feat(455), I2 =>  inp_feat(83), I3 =>  inp_feat(94), I4 =>  inp_feat(289), I5 =>  inp_feat(479), I6 =>  inp_feat(328), I7 =>  inp_feat(494)); 
C_79_S_0_L_6_inst : LUT8 generic map(INIT => "0000010000000000110011000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_0_L_6_out, I0 =>  inp_feat(114), I1 =>  inp_feat(123), I2 =>  inp_feat(359), I3 =>  inp_feat(232), I4 =>  inp_feat(68), I5 =>  inp_feat(270), I6 =>  inp_feat(284), I7 =>  inp_feat(89)); 
C_79_S_0_L_7_inst : LUT8 generic map(INIT => "0000001000000000000000001010000000001000001001000000000000000000000000000000000000000000000100000000000000000000000000000000000010000010100000000000000000000000001010100000101000001010001010100000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_0_L_7_out, I0 =>  inp_feat(94), I1 =>  inp_feat(348), I2 =>  inp_feat(338), I3 =>  inp_feat(469), I4 =>  inp_feat(428), I5 =>  inp_feat(479), I6 =>  inp_feat(420), I7 =>  inp_feat(190)); 
C_79_S_1_L_0_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000001010100000000001100110000000000000011000000000001000000000000000100111000000000") port map( O =>C_79_S_1_L_0_out, I0 =>  inp_feat(23), I1 =>  inp_feat(95), I2 =>  inp_feat(68), I3 =>  inp_feat(141), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_79_S_1_L_1_inst : LUT8 generic map(INIT => "0001000000100000000000000000000000000000000000010000111000000000000000000001000000000000000000000000110100000001000000000000000100000000000000000000000001000100011001000000010100000000000001010000000000000000000000000000000000000001000001010000000100000000") port map( O =>C_79_S_1_L_1_out, I0 =>  inp_feat(479), I1 =>  inp_feat(348), I2 =>  inp_feat(160), I3 =>  inp_feat(474), I4 =>  inp_feat(47), I5 =>  inp_feat(194), I6 =>  inp_feat(451), I7 =>  inp_feat(505)); 
C_79_S_1_L_2_inst : LUT8 generic map(INIT => "1101011100000101000000000000000000000000000001100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_1_L_2_out, I0 =>  inp_feat(79), I1 =>  inp_feat(80), I2 =>  inp_feat(461), I3 =>  inp_feat(16), I4 =>  inp_feat(170), I5 =>  inp_feat(326), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_79_S_1_L_3_inst : LUT8 generic map(INIT => "0000000000000000000000001000000000000000100000001000000010000000000000000000000010000000100000000000000000000000000000000000000000000000100000001000000010000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_1_L_3_out, I0 =>  inp_feat(363), I1 =>  inp_feat(494), I2 =>  inp_feat(128), I3 =>  inp_feat(338), I4 =>  inp_feat(281), I5 =>  inp_feat(171), I6 =>  inp_feat(429), I7 =>  inp_feat(43)); 
C_79_S_1_L_4_inst : LUT8 generic map(INIT => "0000010100000000000000000000000000000111000000000000000100000000000010010000000000000000000000000000110000000000000000000000000010100001000000000000100000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_1_L_4_out, I0 =>  inp_feat(351), I1 =>  inp_feat(160), I2 =>  inp_feat(281), I3 =>  inp_feat(209), I4 =>  inp_feat(89), I5 =>  inp_feat(100), I6 =>  inp_feat(67), I7 =>  inp_feat(25)); 
C_79_S_1_L_5_inst : LUT8 generic map(INIT => "1001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_1_L_5_out, I0 =>  inp_feat(16), I1 =>  inp_feat(294), I2 =>  inp_feat(88), I3 =>  inp_feat(235), I4 =>  inp_feat(501), I5 =>  inp_feat(123), I6 =>  inp_feat(402), I7 =>  inp_feat(303)); 
C_79_S_1_L_6_inst : LUT8 generic map(INIT => "0000000011000000000000000000100010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_1_L_6_out, I0 =>  inp_feat(119), I1 =>  inp_feat(456), I2 =>  inp_feat(207), I3 =>  inp_feat(348), I4 =>  inp_feat(439), I5 =>  inp_feat(47), I6 =>  inp_feat(328), I7 =>  inp_feat(438)); 
C_79_S_1_L_7_inst : LUT8 generic map(INIT => "0000100000000000110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000110000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_1_L_7_out, I0 =>  inp_feat(178), I1 =>  inp_feat(88), I2 =>  inp_feat(256), I3 =>  inp_feat(72), I4 =>  inp_feat(377), I5 =>  inp_feat(13), I6 =>  inp_feat(78), I7 =>  inp_feat(461)); 
C_79_S_2_L_0_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000001010100000000001100110000000000000011000000000001000000000000000100111000000000") port map( O =>C_79_S_2_L_0_out, I0 =>  inp_feat(23), I1 =>  inp_feat(95), I2 =>  inp_feat(68), I3 =>  inp_feat(141), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_79_S_2_L_1_inst : LUT8 generic map(INIT => "0001000000100000000000000000000000000000000000010000111000000000000000000001000000000000000000000000110100000001000000000000000100000000000000000000000001000100011001000000010100000000000001010000000000000000000000000000000000000001000001010000000100000000") port map( O =>C_79_S_2_L_1_out, I0 =>  inp_feat(479), I1 =>  inp_feat(348), I2 =>  inp_feat(160), I3 =>  inp_feat(474), I4 =>  inp_feat(47), I5 =>  inp_feat(194), I6 =>  inp_feat(451), I7 =>  inp_feat(505)); 
C_79_S_2_L_2_inst : LUT8 generic map(INIT => "1000001100101010000000000010001000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_2_L_2_out, I0 =>  inp_feat(27), I1 =>  inp_feat(237), I2 =>  inp_feat(80), I3 =>  inp_feat(461), I4 =>  inp_feat(16), I5 =>  inp_feat(326), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_79_S_2_L_3_inst : LUT8 generic map(INIT => "0001000000011011000000000000100100000000000000000000000000000000000000000010000101000000100001010000000000000000000000000000000000000001001100000100000000000000000000000000000000000000000000000000010000100001000100010000001100000000000000000000000000000000") port map( O =>C_79_S_2_L_3_out, I0 =>  inp_feat(68), I1 =>  inp_feat(479), I2 =>  inp_feat(194), I3 =>  inp_feat(237), I4 =>  inp_feat(502), I5 =>  inp_feat(209), I6 =>  inp_feat(348), I7 =>  inp_feat(43)); 
C_79_S_2_L_4_inst : LUT8 generic map(INIT => "0000010000000000000010101100101000001100000110000000101000001010000000000000000000000000000000000000000010000000000000000000000000000000000010100000000010001000010111000100101000000000000000000000000000000000000010000000000000000000000000000000000000000000") port map( O =>C_79_S_2_L_4_out, I0 =>  inp_feat(67), I1 =>  inp_feat(11), I2 =>  inp_feat(461), I3 =>  inp_feat(348), I4 =>  inp_feat(339), I5 =>  inp_feat(79), I6 =>  inp_feat(121), I7 =>  inp_feat(43)); 
C_79_S_2_L_5_inst : LUT8 generic map(INIT => "0001101100000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000010111000000000000000000000000000010110000000000000000000000000001001100000000000000000000000000000001000000100000000000000000") port map( O =>C_79_S_2_L_5_out, I0 =>  inp_feat(473), I1 =>  inp_feat(281), I2 =>  inp_feat(406), I3 =>  inp_feat(494), I4 =>  inp_feat(399), I5 =>  inp_feat(21), I6 =>  inp_feat(469), I7 =>  inp_feat(81)); 
C_79_S_2_L_6_inst : LUT8 generic map(INIT => "0000000011100000011000001111000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_2_L_6_out, I0 =>  inp_feat(34), I1 =>  inp_feat(206), I2 =>  inp_feat(494), I3 =>  inp_feat(68), I4 =>  inp_feat(237), I5 =>  inp_feat(94), I6 =>  inp_feat(412), I7 =>  inp_feat(98)); 
C_79_S_2_L_7_inst : LUT8 generic map(INIT => "0000000000000000000000000000000011010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000111100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_2_L_7_out, I0 =>  inp_feat(238), I1 =>  inp_feat(485), I2 =>  inp_feat(325), I3 =>  inp_feat(279), I4 =>  inp_feat(400), I5 =>  inp_feat(455), I6 =>  inp_feat(385), I7 =>  inp_feat(80)); 
C_79_S_3_L_0_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000001010100000000001100110000000000000011000000000001000000000000000100111000000000") port map( O =>C_79_S_3_L_0_out, I0 =>  inp_feat(23), I1 =>  inp_feat(95), I2 =>  inp_feat(68), I3 =>  inp_feat(141), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_79_S_3_L_1_inst : LUT8 generic map(INIT => "0010000000000000000000010000100100010000000000000000001000001000000000000000000000001000000000000001000000000000000010110000000100000000000000000000000000000000000000000100010010101111000011010000000000000000000000100000001000000000000000000000101100000010") port map( O =>C_79_S_3_L_1_out, I0 =>  inp_feat(372), I1 =>  inp_feat(348), I2 =>  inp_feat(160), I3 =>  inp_feat(47), I4 =>  inp_feat(194), I5 =>  inp_feat(338), I6 =>  inp_feat(451), I7 =>  inp_feat(505)); 
C_79_S_3_L_2_inst : LUT8 generic map(INIT => "1000001100101010000000000010001000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_3_L_2_out, I0 =>  inp_feat(27), I1 =>  inp_feat(237), I2 =>  inp_feat(80), I3 =>  inp_feat(461), I4 =>  inp_feat(16), I5 =>  inp_feat(326), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_79_S_3_L_3_inst : LUT8 generic map(INIT => "0000000000100000001000001010000000000000000000000000000010000000001010001000000000000000101000000000000000000000000000001000000000000000100000000010000010100000000000001000000000000000000000000000000010000000000000001010000000000000000000000000000010000000") port map( O =>C_79_S_3_L_3_out, I0 =>  inp_feat(415), I1 =>  inp_feat(47), I2 =>  inp_feat(77), I3 =>  inp_feat(455), I4 =>  inp_feat(461), I5 =>  inp_feat(21), I6 =>  inp_feat(469), I7 =>  inp_feat(43)); 
C_79_S_3_L_4_inst : LUT8 generic map(INIT => "1010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_3_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(479), I2 =>  inp_feat(84), I3 =>  inp_feat(136), I4 =>  inp_feat(399), I5 =>  inp_feat(366), I6 =>  inp_feat(72), I7 =>  inp_feat(494)); 
C_79_S_3_L_5_inst : LUT8 generic map(INIT => "0000001000000100000000000000000000000000000000000000000000100000010100100010000000000000000000000000000010000000000000000000000000000000000000110000000000000000000000000000000000000000000000001111001111111111000000000000000000000000000000010000000000000000") port map( O =>C_79_S_3_L_5_out, I0 =>  inp_feat(499), I1 =>  inp_feat(348), I2 =>  inp_feat(97), I3 =>  inp_feat(206), I4 =>  inp_feat(232), I5 =>  inp_feat(95), I6 =>  inp_feat(68), I7 =>  inp_feat(343)); 
C_79_S_3_L_6_inst : LUT8 generic map(INIT => "0000100000000000000000000000000010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_3_L_6_out, I0 =>  inp_feat(420), I1 =>  inp_feat(422), I2 =>  inp_feat(348), I3 =>  inp_feat(280), I4 =>  inp_feat(147), I5 =>  inp_feat(281), I6 =>  inp_feat(123), I7 =>  inp_feat(406)); 
C_79_S_3_L_7_inst : LUT8 generic map(INIT => "0001000000000000000101000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011000000100000000000000010000000000000000000000000000000000000001100000001000000000000001000000000000000000000000000000000000000") port map( O =>C_79_S_3_L_7_out, I0 =>  inp_feat(160), I1 =>  inp_feat(388), I2 =>  inp_feat(102), I3 =>  inp_feat(290), I4 =>  inp_feat(429), I5 =>  inp_feat(164), I6 =>  inp_feat(438), I7 =>  inp_feat(338)); 
C_79_S_4_L_0_inst : LUT8 generic map(INIT => "0000010000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000001010100000000001100110000000000000011000000000001000000000000000100111000000000") port map( O =>C_79_S_4_L_0_out, I0 =>  inp_feat(23), I1 =>  inp_feat(95), I2 =>  inp_feat(68), I3 =>  inp_feat(141), I4 =>  inp_feat(160), I5 =>  inp_feat(206), I6 =>  inp_feat(479), I7 =>  inp_feat(237)); 
C_79_S_4_L_1_inst : LUT8 generic map(INIT => "0010000000000000000000010000100100010000000000000000001000001000000000000000000000001000000000000001000000000000000010110000000100000000000000000000000000000000000000000100010010101111000011010000000000000000000000100000001000000000000000000000101100000010") port map( O =>C_79_S_4_L_1_out, I0 =>  inp_feat(372), I1 =>  inp_feat(348), I2 =>  inp_feat(160), I3 =>  inp_feat(47), I4 =>  inp_feat(194), I5 =>  inp_feat(338), I6 =>  inp_feat(451), I7 =>  inp_feat(505)); 
C_79_S_4_L_2_inst : LUT8 generic map(INIT => "1000001100101010000000000010001000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_4_L_2_out, I0 =>  inp_feat(27), I1 =>  inp_feat(237), I2 =>  inp_feat(80), I3 =>  inp_feat(461), I4 =>  inp_feat(16), I5 =>  inp_feat(326), I6 =>  inp_feat(283), I7 =>  inp_feat(494)); 
C_79_S_4_L_3_inst : LUT8 generic map(INIT => "0000000000100000001000001010000000000000000000000000000010000000001010001000000000000000101000000000000000000000000000001000000000000000100000000010000010100000000000001000000000000000000000000000000010000000000000001010000000000000000000000000000010000000") port map( O =>C_79_S_4_L_3_out, I0 =>  inp_feat(415), I1 =>  inp_feat(47), I2 =>  inp_feat(77), I3 =>  inp_feat(455), I4 =>  inp_feat(461), I5 =>  inp_feat(21), I6 =>  inp_feat(469), I7 =>  inp_feat(43)); 
C_79_S_4_L_4_inst : LUT8 generic map(INIT => "1010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_4_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(479), I2 =>  inp_feat(84), I3 =>  inp_feat(136), I4 =>  inp_feat(399), I5 =>  inp_feat(366), I6 =>  inp_feat(72), I7 =>  inp_feat(494)); 
C_79_S_4_L_5_inst : LUT8 generic map(INIT => "0110000000000001000000000000000000000000000000001100000000010000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000001111000011000000001000000000000001000000000000000000000001000000111100000000000000000000") port map( O =>C_79_S_4_L_5_out, I0 =>  inp_feat(348), I1 =>  inp_feat(295), I2 =>  inp_feat(487), I3 =>  inp_feat(265), I4 =>  inp_feat(67), I5 =>  inp_feat(68), I6 =>  inp_feat(261), I7 =>  inp_feat(343)); 
C_79_S_4_L_6_inst : LUT8 generic map(INIT => "0000001000000000100100001001000100000000001000000000000000000000010101110000110101110001001011110000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") port map( O =>C_79_S_4_L_6_out, I0 =>  inp_feat(248), I1 =>  inp_feat(348), I2 =>  inp_feat(25), I3 =>  inp_feat(206), I4 =>  inp_feat(6), I5 =>  inp_feat(232), I6 =>  inp_feat(338), I7 =>  inp_feat(375)); 
C_79_S_4_L_7_inst : LUT8 generic map(INIT => "0110000000001000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010110000011110000001000000010000100100001111001100010000001100110000000000000000000000000000000000000001000000000000000000000000") port map( O =>C_79_S_4_L_7_out, I0 =>  inp_feat(348), I1 =>  inp_feat(80), I2 =>  inp_feat(365), I3 =>  inp_feat(338), I4 =>  inp_feat(319), I5 =>  inp_feat(100), I6 =>  inp_feat(102), I7 =>  inp_feat(281)); 

C_0_S_0_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_0_S_0_out, I0 =>  C_0_S_0_L_0_out, I1 =>  C_0_S_0_L_1_out, I2 =>  C_0_S_0_L_2_out, I3 =>  C_0_S_0_L_3_out, I4 =>  C_0_S_0_L_4_out, I5 =>  C_0_S_0_L_5_out, I6 =>  C_0_S_0_L_6_out, I7 =>  C_0_S_0_L_7_out); 
C_0_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000000000000") port map( O =>C_0_S_1_out, I0 =>  C_0_S_1_L_0_out, I1 =>  C_0_S_1_L_1_out, I2 =>  C_0_S_1_L_2_out, I3 =>  C_0_S_1_L_3_out, I4 =>  C_0_S_1_L_4_out, I5 =>  C_0_S_1_L_5_out, I6 =>  C_0_S_1_L_6_out, I7 =>  C_0_S_1_L_7_out); 
C_0_S_2_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_0_S_2_out, I0 =>  C_0_S_2_L_0_out, I1 =>  C_0_S_2_L_1_out, I2 =>  C_0_S_2_L_2_out, I3 =>  C_0_S_2_L_3_out, I4 =>  C_0_S_2_L_4_out, I5 =>  C_0_S_2_L_5_out, I6 =>  C_0_S_2_L_6_out, I7 =>  C_0_S_2_L_7_out); 
C_0_S_3_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_0_S_3_out, I0 =>  C_0_S_3_L_0_out, I1 =>  C_0_S_3_L_1_out, I2 =>  C_0_S_3_L_2_out, I3 =>  C_0_S_3_L_3_out, I4 =>  C_0_S_3_L_4_out, I5 =>  C_0_S_3_L_5_out, I6 =>  C_0_S_3_L_6_out, I7 =>  C_0_S_3_L_7_out); 
C_0_S_4_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_0_S_4_out, I0 =>  C_0_S_4_L_0_out, I1 =>  C_0_S_4_L_1_out, I2 =>  C_0_S_4_L_2_out, I3 =>  C_0_S_4_L_3_out, I4 =>  C_0_S_4_L_4_out, I5 =>  C_0_S_4_L_5_out, I6 =>  C_0_S_4_L_6_out, I7 =>  C_0_S_4_L_7_out); 

C_0_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_0_out, I0 =>  C_0_S_0_out, I1 =>  C_0_S_1_out, I2 =>  C_0_S_2_out, I3 =>  C_0_S_3_out, I4 =>  C_0_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_1_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111010101110101010101000111111101110111011101010111010001110101010101000101010001000000011111110111010101110101010101000111010001010100010001000100000001110101010101000101010001000000010001000100000001000000000000000") port map( O =>C_1_S_0_out, I0 =>  C_1_S_0_L_0_out, I1 =>  C_1_S_0_L_1_out, I2 =>  C_1_S_0_L_2_out, I3 =>  C_1_S_0_L_3_out, I4 =>  C_1_S_0_L_4_out, I5 =>  C_1_S_0_L_5_out, I6 =>  C_1_S_0_L_6_out, I7 =>  C_1_S_0_L_7_out); 
C_1_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111011101110101011101010100010001110100010001000100010001000000011111110111011101110111011101000111011101010100010101000100010001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_1_S_1_out, I0 =>  C_1_S_1_L_0_out, I1 =>  C_1_S_1_L_1_out, I2 =>  C_1_S_1_L_2_out, I3 =>  C_1_S_1_L_3_out, I4 =>  C_1_S_1_L_4_out, I5 =>  C_1_S_1_L_5_out, I6 =>  C_1_S_1_L_6_out, I7 =>  C_1_S_1_L_7_out); 
C_1_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011101110111010101110101010101000111011101110101011101010101010001110100010001000100010001000000011111110111011101110111011101000111010101010100010101000100010001110101010101000101010001000100010101000100000001000000000000000") port map( O =>C_1_S_2_out, I0 =>  C_1_S_2_L_0_out, I1 =>  C_1_S_2_L_1_out, I2 =>  C_1_S_2_L_2_out, I3 =>  C_1_S_2_L_3_out, I4 =>  C_1_S_2_L_4_out, I5 =>  C_1_S_2_L_5_out, I6 =>  C_1_S_2_L_6_out, I7 =>  C_1_S_2_L_7_out); 
C_1_S_3_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111011101110100011101000101010001110100010001000100010001000000011111110111011101110111011101000111010101110100011101000100010001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_1_S_3_out, I0 =>  C_1_S_3_L_0_out, I1 =>  C_1_S_3_L_1_out, I2 =>  C_1_S_3_L_2_out, I3 =>  C_1_S_3_L_3_out, I4 =>  C_1_S_3_L_4_out, I5 =>  C_1_S_3_L_5_out, I6 =>  C_1_S_3_L_6_out, I7 =>  C_1_S_3_L_7_out); 
C_1_S_4_inst : LUT8 generic map(INIT => "1111111011111110111011101110101011101110111010101110100010101000111011101110101011101000101010001110100010101000100010001000000011111110111011101110101011101000111010101110100010101000100010001110101011101000101010001000100010101000100010001000000010000000") port map( O =>C_1_S_4_out, I0 =>  C_1_S_4_L_0_out, I1 =>  C_1_S_4_L_1_out, I2 =>  C_1_S_4_L_2_out, I3 =>  C_1_S_4_L_3_out, I4 =>  C_1_S_4_L_4_out, I5 =>  C_1_S_4_L_5_out, I6 =>  C_1_S_4_L_6_out, I7 =>  C_1_S_4_L_7_out); 

C_1_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_1_out, I0 =>  C_1_S_0_out, I1 =>  C_1_S_1_out, I2 =>  C_1_S_2_out, I3 =>  C_1_S_3_out, I4 =>  C_1_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_2_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111111111110001111100010000000111111111111100011111000100000001111111011101000111010001000000011111110111010001110100010000000111111101110000011100000000000001111111011100000111000000000000011101000100000001000000000000000") port map( O =>C_2_S_0_out, I0 =>  C_2_S_0_L_0_out, I1 =>  C_2_S_0_L_1_out, I2 =>  C_2_S_0_L_2_out, I3 =>  C_2_S_0_L_3_out, I4 =>  C_2_S_0_L_4_out, I5 =>  C_2_S_0_L_5_out, I6 =>  C_2_S_0_L_6_out, I7 =>  C_2_S_0_L_7_out); 
C_2_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001111100010100000111111101110100011111000101000001111101011100000111010001000000011111110111010001111100010100000111110101110000011101000100000001111101011100000111010001000000011101000100000001000000000000000") port map( O =>C_2_S_1_out, I0 =>  C_2_S_1_L_0_out, I1 =>  C_2_S_1_L_1_out, I2 =>  C_2_S_1_L_2_out, I3 =>  C_2_S_1_L_3_out, I4 =>  C_2_S_1_L_4_out, I5 =>  C_2_S_1_L_5_out, I6 =>  C_2_S_1_L_6_out, I7 =>  C_2_S_1_L_7_out); 
C_2_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010100000111111101110100011101000100000001111101011101000111010001000000011111110111010001110100010100000111111101110100011101000100000001111101011101000111010001000000011101000100000001000000000000000") port map( O =>C_2_S_2_out, I0 =>  C_2_S_2_L_0_out, I1 =>  C_2_S_2_L_1_out, I2 =>  C_2_S_2_L_2_out, I3 =>  C_2_S_2_L_3_out, I4 =>  C_2_S_2_L_4_out, I5 =>  C_2_S_2_L_5_out, I6 =>  C_2_S_2_L_6_out, I7 =>  C_2_S_2_L_7_out); 
C_2_S_3_inst : LUT8 generic map(INIT => "1111111111111010111111101110100011111110111010001111101010100000111111101110100011111010101000001111101010100000111010001000000011111110111010001111101010100000111110101010000011101000100000001111101010100000111010001000000011101000100000001010000000000000") port map( O =>C_2_S_3_out, I0 =>  C_2_S_3_L_0_out, I1 =>  C_2_S_3_L_1_out, I2 =>  C_2_S_3_L_2_out, I3 =>  C_2_S_3_L_3_out, I4 =>  C_2_S_3_L_4_out, I5 =>  C_2_S_3_L_5_out, I6 =>  C_2_S_3_L_6_out, I7 =>  C_2_S_3_L_7_out); 
C_2_S_4_inst : LUT8 generic map(INIT => "1111111111111110111110101110100011111110111110101110100010100000111111101111100011101000100000001111111011101000111000001000000011111110111110001110100010000000111111101110100011100000100000001111101011101000101000001000000011101000101000001000000000000000") port map( O =>C_2_S_4_out, I0 =>  C_2_S_4_L_0_out, I1 =>  C_2_S_4_L_1_out, I2 =>  C_2_S_4_L_2_out, I3 =>  C_2_S_4_L_3_out, I4 =>  C_2_S_4_L_4_out, I5 =>  C_2_S_4_L_5_out, I6 =>  C_2_S_4_L_6_out, I7 =>  C_2_S_4_L_7_out); 

C_2_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_2_out, I0 =>  C_2_S_0_out, I1 =>  C_2_S_1_out, I2 =>  C_2_S_2_out, I3 =>  C_2_S_3_out, I4 =>  C_2_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_3_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101110101010101110101010101000111010101010101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101010101010001110101010101000101010101000100010101010101010001010100010001000") port map( O =>C_3_S_0_out, I0 =>  C_3_S_0_L_0_out, I1 =>  C_3_S_0_L_1_out, I2 =>  C_3_S_0_L_2_out, I3 =>  C_3_S_0_L_3_out, I4 =>  C_3_S_0_L_4_out, I5 =>  C_3_S_0_L_5_out, I6 =>  C_3_S_0_L_6_out, I7 =>  C_3_S_0_L_7_out); 
C_3_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_3_S_1_out, I0 =>  C_3_S_1_L_0_out, I1 =>  C_3_S_1_L_1_out, I2 =>  C_3_S_1_L_2_out, I3 =>  C_3_S_1_L_3_out, I4 =>  C_3_S_1_L_4_out, I5 =>  C_3_S_1_L_5_out, I6 =>  C_3_S_1_L_6_out, I7 =>  C_3_S_1_L_7_out); 
C_3_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001000000010001000100000001000000000000000") port map( O =>C_3_S_2_out, I0 =>  C_3_S_2_L_0_out, I1 =>  C_3_S_2_L_1_out, I2 =>  C_3_S_2_L_2_out, I3 =>  C_3_S_2_L_3_out, I4 =>  C_3_S_2_L_4_out, I5 =>  C_3_S_2_L_5_out, I6 =>  C_3_S_2_L_6_out, I7 =>  C_3_S_2_L_7_out); 
C_3_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101110110011001000111111111111110011101100110010001110110011001000110000000000000011111111111111001110110011001000111011001100100011000000000000001110110011001000100000000000000010000000000000000000000000000000") port map( O =>C_3_S_3_out, I0 =>  C_3_S_3_L_0_out, I1 =>  C_3_S_3_L_1_out, I2 =>  C_3_S_3_L_2_out, I3 =>  C_3_S_3_L_3_out, I4 =>  C_3_S_3_L_4_out, I5 =>  C_3_S_3_L_5_out, I6 =>  C_3_S_3_L_6_out, I7 =>  C_3_S_3_L_7_out); 
C_3_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011101110111010001110110011101000111111101110111011101110111010001110100011001000111010001000100011101110111010001110110011101000111010001000100010001000100000001110100011001000111010001000100010001000100000001000000000000000") port map( O =>C_3_S_4_out, I0 =>  C_3_S_4_L_0_out, I1 =>  C_3_S_4_L_1_out, I2 =>  C_3_S_4_L_2_out, I3 =>  C_3_S_4_L_3_out, I4 =>  C_3_S_4_L_4_out, I5 =>  C_3_S_4_L_5_out, I6 =>  C_3_S_4_L_6_out, I7 =>  C_3_S_4_L_7_out); 

C_3_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_3_out, I0 =>  C_3_S_0_out, I1 =>  C_3_S_1_out, I2 =>  C_3_S_2_out, I3 =>  C_3_S_3_out, I4 =>  C_3_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_4_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101110101011101010111010101110101010101000111010101110101011101010101010001110101010101000101010001010100011101010111010101110101010101000111010101010100010101000101010001110101010101000101010001010100010101000101010001010100010001000") port map( O =>C_4_S_0_out, I0 =>  C_4_S_0_L_0_out, I1 =>  C_4_S_0_L_1_out, I2 =>  C_4_S_0_L_2_out, I3 =>  C_4_S_0_L_3_out, I4 =>  C_4_S_0_L_4_out, I5 =>  C_4_S_0_L_5_out, I6 =>  C_4_S_0_L_6_out, I7 =>  C_4_S_0_L_7_out); 
C_4_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110101011101110101010001110101010101000111010001000000011111110111010001110101010101000111010101000100010101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_4_S_1_out, I0 =>  C_4_S_1_L_0_out, I1 =>  C_4_S_1_L_1_out, I2 =>  C_4_S_1_L_2_out, I3 =>  C_4_S_1_L_3_out, I4 =>  C_4_S_1_L_4_out, I5 =>  C_4_S_1_L_5_out, I6 =>  C_4_S_1_L_6_out, I7 =>  C_4_S_1_L_7_out); 
C_4_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110110011111110111011001110100011001000111111101110111011101100111010001110110011101000110010001000000011111110111011001110100011001000111010001100100010001000100000001110110011101000110010001000000011001000100000001000000000000000") port map( O =>C_4_S_2_out, I0 =>  C_4_S_2_L_0_out, I1 =>  C_4_S_2_L_1_out, I2 =>  C_4_S_2_L_2_out, I3 =>  C_4_S_2_L_3_out, I4 =>  C_4_S_2_L_4_out, I5 =>  C_4_S_2_L_5_out, I6 =>  C_4_S_2_L_6_out, I7 =>  C_4_S_2_L_7_out); 
C_4_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110100010001000111111101110101011101000101010001110100010101000100010001000000011111110111011101110101011101000111010101110100010101000100000001110111011101000101010001000000010101000100000001000000000000000") port map( O =>C_4_S_3_out, I0 =>  C_4_S_3_L_0_out, I1 =>  C_4_S_3_L_1_out, I2 =>  C_4_S_3_L_2_out, I3 =>  C_4_S_3_L_3_out, I4 =>  C_4_S_3_L_4_out, I5 =>  C_4_S_3_L_5_out, I6 =>  C_4_S_3_L_6_out, I7 =>  C_4_S_3_L_7_out); 
C_4_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111101110100011111111111110101110100010000000111111111111111011111010101000001111111011100000101000000000000011111111111110101111100010000000111110101010000010000000000000001111111011101000101000000000000011101000100000000000000000000000") port map( O =>C_4_S_4_out, I0 =>  C_4_S_4_L_0_out, I1 =>  C_4_S_4_L_1_out, I2 =>  C_4_S_4_L_2_out, I3 =>  C_4_S_4_L_3_out, I4 =>  C_4_S_4_L_4_out, I5 =>  C_4_S_4_L_5_out, I6 =>  C_4_S_4_L_6_out, I7 =>  C_4_S_4_L_7_out); 

C_4_inst : LUT8 generic map(INIT => "1110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000") port map( O =>C_4_out, I0 =>  C_4_S_0_out, I1 =>  C_4_S_1_out, I2 =>  C_4_S_2_out, I3 =>  C_4_S_3_out, I4 =>  C_4_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_5_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101000111010101110101011101010101010001110101010101000101010001010100011101010111010101110101010101000111010101010100010101000101010001110101010101010101010101010100010101010101010001010100010000000") port map( O =>C_5_S_0_out, I0 =>  C_5_S_0_L_0_out, I1 =>  C_5_S_0_L_1_out, I2 =>  C_5_S_0_L_2_out, I3 =>  C_5_S_0_L_3_out, I4 =>  C_5_S_0_L_4_out, I5 =>  C_5_S_0_L_5_out, I6 =>  C_5_S_0_L_6_out, I7 =>  C_5_S_0_L_7_out); 
C_5_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011111110101010001111111010101000111010001000000011111110111010001110101010000000111010101000000011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_5_S_1_out, I0 =>  C_5_S_1_L_0_out, I1 =>  C_5_S_1_L_1_out, I2 =>  C_5_S_1_L_2_out, I3 =>  C_5_S_1_L_3_out, I4 =>  C_5_S_1_L_4_out, I5 =>  C_5_S_1_L_5_out, I6 =>  C_5_S_1_L_6_out, I7 =>  C_5_S_1_L_7_out); 
C_5_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111101111100011111110111111101111100011100000111111101111100011101000110000001111100011100000100000001000000011111110111111101111100011100000111111001110100011100000100000001111100011100000100000001000000011100000100000000000000000000000") port map( O =>C_5_S_2_out, I0 =>  C_5_S_2_L_0_out, I1 =>  C_5_S_2_L_1_out, I2 =>  C_5_S_2_L_2_out, I3 =>  C_5_S_2_L_3_out, I4 =>  C_5_S_2_L_4_out, I5 =>  C_5_S_2_L_5_out, I6 =>  C_5_S_2_L_6_out, I7 =>  C_5_S_2_L_7_out); 
C_5_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111110101011111111111011101110101010000000111111111110111011101110100010001110111010001000100010000000000011111111111011101110111010001000111011101000100010001000000000001111111010101000100010000000000010101000000000000000000000000000") port map( O =>C_5_S_3_out, I0 =>  C_5_S_3_L_0_out, I1 =>  C_5_S_3_L_1_out, I2 =>  C_5_S_3_L_2_out, I3 =>  C_5_S_3_L_3_out, I4 =>  C_5_S_3_L_4_out, I5 =>  C_5_S_3_L_5_out, I6 =>  C_5_S_3_L_6_out, I7 =>  C_5_S_3_L_7_out); 
C_5_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111101111111011111110111010101110100010000000111111111111111011101010101010001110100010000000100000000000000011111111111111101111111011101000111010101010100010000000000000001111111011101000101010001000000010000000100000000000000000000000") port map( O =>C_5_S_4_out, I0 =>  C_5_S_4_L_0_out, I1 =>  C_5_S_4_L_1_out, I2 =>  C_5_S_4_L_2_out, I3 =>  C_5_S_4_L_3_out, I4 =>  C_5_S_4_L_4_out, I5 =>  C_5_S_4_L_5_out, I6 =>  C_5_S_4_L_6_out, I7 =>  C_5_S_4_L_7_out); 

C_5_inst : LUT8 generic map(INIT => "1110111010101000111010101000100011101110101010001110101010001000111011101010100011101010100010001110111010101000111010101000100011101110101010001110101010001000111011101010100011101010100010001110111010101000111010101000100011101110101010001110101010001000") port map( O =>C_5_out, I0 =>  C_5_S_0_out, I1 =>  C_5_S_1_out, I2 =>  C_5_S_2_out, I3 =>  C_5_S_3_out, I4 =>  C_5_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_6_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_6_S_0_out, I0 =>  C_6_S_0_L_0_out, I1 =>  C_6_S_0_L_1_out, I2 =>  C_6_S_0_L_2_out, I3 =>  C_6_S_0_L_3_out, I4 =>  C_6_S_0_L_4_out, I5 =>  C_6_S_0_L_5_out, I6 =>  C_6_S_0_L_6_out, I7 =>  C_6_S_0_L_7_out); 
C_6_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_6_S_1_out, I0 =>  C_6_S_1_L_0_out, I1 =>  C_6_S_1_L_1_out, I2 =>  C_6_S_1_L_2_out, I3 =>  C_6_S_1_L_3_out, I4 =>  C_6_S_1_L_4_out, I5 =>  C_6_S_1_L_5_out, I6 =>  C_6_S_1_L_6_out, I7 =>  C_6_S_1_L_7_out); 
C_6_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_6_S_2_out, I0 =>  C_6_S_2_L_0_out, I1 =>  C_6_S_2_L_1_out, I2 =>  C_6_S_2_L_2_out, I3 =>  C_6_S_2_L_3_out, I4 =>  C_6_S_2_L_4_out, I5 =>  C_6_S_2_L_5_out, I6 =>  C_6_S_2_L_6_out, I7 =>  C_6_S_2_L_7_out); 
C_6_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_6_S_3_out, I0 =>  C_6_S_3_L_0_out, I1 =>  C_6_S_3_L_1_out, I2 =>  C_6_S_3_L_2_out, I3 =>  C_6_S_3_L_3_out, I4 =>  C_6_S_3_L_4_out, I5 =>  C_6_S_3_L_5_out, I6 =>  C_6_S_3_L_6_out, I7 =>  C_6_S_3_L_7_out); 
C_6_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_6_S_4_out, I0 =>  C_6_S_4_L_0_out, I1 =>  C_6_S_4_L_1_out, I2 =>  C_6_S_4_L_2_out, I3 =>  C_6_S_4_L_3_out, I4 =>  C_6_S_4_L_4_out, I5 =>  C_6_S_4_L_5_out, I6 =>  C_6_S_4_L_6_out, I7 =>  C_6_S_4_L_7_out); 

C_6_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_6_out, I0 =>  C_6_S_0_out, I1 =>  C_6_S_1_out, I2 =>  C_6_S_2_out, I3 =>  C_6_S_3_out, I4 =>  C_6_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_7_S_0_inst : LUT8 generic map(INIT => "1110111011101110111011101010100011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100011101010100010001000100010001000") port map( O =>C_7_S_0_out, I0 =>  C_7_S_0_L_0_out, I1 =>  C_7_S_0_L_1_out, I2 =>  C_7_S_0_L_2_out, I3 =>  C_7_S_0_L_3_out, I4 =>  C_7_S_0_L_4_out, I5 =>  C_7_S_0_L_5_out, I6 =>  C_7_S_0_L_6_out, I7 =>  C_7_S_0_L_7_out); 
C_7_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001111101010000000111111101110100011111010100000001111101010000000111010000000000011111111111010001111111010100000111111101010000011101000100000001111111010100000111010001000000011101000100000001000000000000000") port map( O =>C_7_S_1_out, I0 =>  C_7_S_1_L_0_out, I1 =>  C_7_S_1_L_1_out, I2 =>  C_7_S_1_L_2_out, I3 =>  C_7_S_1_L_3_out, I4 =>  C_7_S_1_L_4_out, I5 =>  C_7_S_1_L_5_out, I6 =>  C_7_S_1_L_6_out, I7 =>  C_7_S_1_L_7_out); 
C_7_S_2_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100010101000111111101110100011101000101010001110101010101000101010001000000011111110111010101110101010101000111010101110100011101000100000001110101011101000111010001000000011101000100000001000000010000000") port map( O =>C_7_S_2_out, I0 =>  C_7_S_2_L_0_out, I1 =>  C_7_S_2_L_1_out, I2 =>  C_7_S_2_L_2_out, I3 =>  C_7_S_2_L_3_out, I4 =>  C_7_S_2_L_4_out, I5 =>  C_7_S_2_L_5_out, I6 =>  C_7_S_2_L_6_out, I7 =>  C_7_S_2_L_7_out); 
C_7_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111111111100011111111111110001111111010100000111111111111101011111110111000001111111111100000111110000000000011111111111000001111100000000000111110001000000010100000000000001111101010000000111000000000000011100000000000001000000000000000") port map( O =>C_7_S_3_out, I0 =>  C_7_S_3_L_0_out, I1 =>  C_7_S_3_L_1_out, I2 =>  C_7_S_3_L_2_out, I3 =>  C_7_S_3_L_3_out, I4 =>  C_7_S_3_L_4_out, I5 =>  C_7_S_3_L_5_out, I6 =>  C_7_S_3_L_6_out, I7 =>  C_7_S_3_L_7_out); 
C_7_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101111110011111110111111001111110011101000111111001110100011101000110000001110100011000000110010001000000011111110111011001111110011101000111111001110100011101000110000001110100011000000110000001000000011000000100000001000000000000000") port map( O =>C_7_S_4_out, I0 =>  C_7_S_4_L_0_out, I1 =>  C_7_S_4_L_1_out, I2 =>  C_7_S_4_L_2_out, I3 =>  C_7_S_4_L_3_out, I4 =>  C_7_S_4_L_4_out, I5 =>  C_7_S_4_L_5_out, I6 =>  C_7_S_4_L_6_out, I7 =>  C_7_S_4_L_7_out); 

C_7_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_7_out, I0 =>  C_7_S_0_out, I1 =>  C_7_S_1_out, I2 =>  C_7_S_2_out, I3 =>  C_7_S_3_out, I4 =>  C_7_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_8_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_8_S_0_out, I0 =>  C_8_S_0_L_0_out, I1 =>  C_8_S_0_L_1_out, I2 =>  C_8_S_0_L_2_out, I3 =>  C_8_S_0_L_3_out, I4 =>  C_8_S_0_L_4_out, I5 =>  C_8_S_0_L_5_out, I6 =>  C_8_S_0_L_6_out, I7 =>  C_8_S_0_L_7_out); 
C_8_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_8_S_1_out, I0 =>  C_8_S_1_L_0_out, I1 =>  C_8_S_1_L_1_out, I2 =>  C_8_S_1_L_2_out, I3 =>  C_8_S_1_L_3_out, I4 =>  C_8_S_1_L_4_out, I5 =>  C_8_S_1_L_5_out, I6 =>  C_8_S_1_L_6_out, I7 =>  C_8_S_1_L_7_out); 
C_8_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_8_S_2_out, I0 =>  C_8_S_2_L_0_out, I1 =>  C_8_S_2_L_1_out, I2 =>  C_8_S_2_L_2_out, I3 =>  C_8_S_2_L_3_out, I4 =>  C_8_S_2_L_4_out, I5 =>  C_8_S_2_L_5_out, I6 =>  C_8_S_2_L_6_out, I7 =>  C_8_S_2_L_7_out); 
C_8_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_8_S_3_out, I0 =>  C_8_S_3_L_0_out, I1 =>  C_8_S_3_L_1_out, I2 =>  C_8_S_3_L_2_out, I3 =>  C_8_S_3_L_3_out, I4 =>  C_8_S_3_L_4_out, I5 =>  C_8_S_3_L_5_out, I6 =>  C_8_S_3_L_6_out, I7 =>  C_8_S_3_L_7_out); 
C_8_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_8_S_4_out, I0 =>  C_8_S_4_L_0_out, I1 =>  C_8_S_4_L_1_out, I2 =>  C_8_S_4_L_2_out, I3 =>  C_8_S_4_L_3_out, I4 =>  C_8_S_4_L_4_out, I5 =>  C_8_S_4_L_5_out, I6 =>  C_8_S_4_L_6_out, I7 =>  C_8_S_4_L_7_out); 

C_8_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_8_out, I0 =>  C_8_S_0_out, I1 =>  C_8_S_1_out, I2 =>  C_8_S_2_out, I3 =>  C_8_S_3_out, I4 =>  C_8_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_9_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_9_S_0_out, I0 =>  C_9_S_0_L_0_out, I1 =>  C_9_S_0_L_1_out, I2 =>  C_9_S_0_L_2_out, I3 =>  C_9_S_0_L_3_out, I4 =>  C_9_S_0_L_4_out, I5 =>  C_9_S_0_L_5_out, I6 =>  C_9_S_0_L_6_out, I7 =>  C_9_S_0_L_7_out); 
C_9_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_9_S_1_out, I0 =>  C_9_S_1_L_0_out, I1 =>  C_9_S_1_L_1_out, I2 =>  C_9_S_1_L_2_out, I3 =>  C_9_S_1_L_3_out, I4 =>  C_9_S_1_L_4_out, I5 =>  C_9_S_1_L_5_out, I6 =>  C_9_S_1_L_6_out, I7 =>  C_9_S_1_L_7_out); 
C_9_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_9_S_2_out, I0 =>  C_9_S_2_L_0_out, I1 =>  C_9_S_2_L_1_out, I2 =>  C_9_S_2_L_2_out, I3 =>  C_9_S_2_L_3_out, I4 =>  C_9_S_2_L_4_out, I5 =>  C_9_S_2_L_5_out, I6 =>  C_9_S_2_L_6_out, I7 =>  C_9_S_2_L_7_out); 
C_9_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_9_S_3_out, I0 =>  C_9_S_3_L_0_out, I1 =>  C_9_S_3_L_1_out, I2 =>  C_9_S_3_L_2_out, I3 =>  C_9_S_3_L_3_out, I4 =>  C_9_S_3_L_4_out, I5 =>  C_9_S_3_L_5_out, I6 =>  C_9_S_3_L_6_out, I7 =>  C_9_S_3_L_7_out); 
C_9_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_9_S_4_out, I0 =>  C_9_S_4_L_0_out, I1 =>  C_9_S_4_L_1_out, I2 =>  C_9_S_4_L_2_out, I3 =>  C_9_S_4_L_3_out, I4 =>  C_9_S_4_L_4_out, I5 =>  C_9_S_4_L_5_out, I6 =>  C_9_S_4_L_6_out, I7 =>  C_9_S_4_L_7_out); 

C_9_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_9_out, I0 =>  C_9_S_0_out, I1 =>  C_9_S_1_out, I2 =>  C_9_S_2_out, I3 =>  C_9_S_3_out, I4 =>  C_9_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_10_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101110100011101010111010101110101010101000111010101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000101010001110101010101000101010001010100011101000101010001010100010000000") port map( O =>C_10_S_0_out, I0 =>  C_10_S_0_L_0_out, I1 =>  C_10_S_0_L_1_out, I2 =>  C_10_S_0_L_2_out, I3 =>  C_10_S_0_L_3_out, I4 =>  C_10_S_0_L_4_out, I5 =>  C_10_S_0_L_5_out, I6 =>  C_10_S_0_L_6_out, I7 =>  C_10_S_0_L_7_out); 
C_10_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101000111111101110101010101010101010101010101010101000101010001000000011111110111010101110101010101010101010101010101010101000100000001110101010101010101010101010100010101010101010001010100010000000") port map( O =>C_10_S_1_out, I0 =>  C_10_S_1_L_0_out, I1 =>  C_10_S_1_L_1_out, I2 =>  C_10_S_1_L_2_out, I3 =>  C_10_S_1_L_3_out, I4 =>  C_10_S_1_L_4_out, I5 =>  C_10_S_1_L_5_out, I6 =>  C_10_S_1_L_6_out, I7 =>  C_10_S_1_L_7_out); 
C_10_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111101111100011111110111110001111100011100000111111101111110011111000111000001111100011100000110000000000000011111111111111001111100011100000111110001110000011000000100000001111100011100000111000001000000011100000100000000000000000000000") port map( O =>C_10_S_2_out, I0 =>  C_10_S_2_L_0_out, I1 =>  C_10_S_2_L_1_out, I2 =>  C_10_S_2_L_2_out, I3 =>  C_10_S_2_L_3_out, I4 =>  C_10_S_2_L_4_out, I5 =>  C_10_S_2_L_5_out, I6 =>  C_10_S_2_L_6_out, I7 =>  C_10_S_2_L_7_out); 
C_10_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010101110100010000000111111101110100011101000100000001110101010001000100000000000000011111111111111101110111010101000111111101110100011101000100000001111111011101000101010001000000011101000100000001000000000000000") port map( O =>C_10_S_3_out, I0 =>  C_10_S_3_L_0_out, I1 =>  C_10_S_3_L_1_out, I2 =>  C_10_S_3_L_2_out, I3 =>  C_10_S_3_L_3_out, I4 =>  C_10_S_3_L_4_out, I5 =>  C_10_S_3_L_5_out, I6 =>  C_10_S_3_L_6_out, I7 =>  C_10_S_3_L_7_out); 
C_10_S_4_inst : LUT8 generic map(INIT => "1111111011111110111111101110101011111010111010101110101011101000111110101110100011101000101010001110100010101000101010001000000011111110111010101110101011101000111010101110100011101000101000001110100010101000101010001010000010101000100000001000000010000000") port map( O =>C_10_S_4_out, I0 =>  C_10_S_4_L_0_out, I1 =>  C_10_S_4_L_1_out, I2 =>  C_10_S_4_L_2_out, I3 =>  C_10_S_4_L_3_out, I4 =>  C_10_S_4_L_4_out, I5 =>  C_10_S_4_L_5_out, I6 =>  C_10_S_4_L_6_out, I7 =>  C_10_S_4_L_7_out); 

C_10_inst : LUT8 generic map(INIT => "1110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000") port map( O =>C_10_out, I0 =>  C_10_S_0_out, I1 =>  C_10_S_1_out, I2 =>  C_10_S_2_out, I3 =>  C_10_S_3_out, I4 =>  C_10_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_11_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101110100010001000111111111111111011101100110010001111111011101000100000000000000011111111111111101110100010000000111011001100100010000000000000001110111011101000100000000000000010000000000000000000000000000000") port map( O =>C_11_S_0_out, I0 =>  C_11_S_0_L_0_out, I1 =>  C_11_S_0_L_1_out, I2 =>  C_11_S_0_L_2_out, I3 =>  C_11_S_0_L_3_out, I4 =>  C_11_S_0_L_4_out, I5 =>  C_11_S_0_L_5_out, I6 =>  C_11_S_0_L_6_out, I7 =>  C_11_S_0_L_7_out); 
C_11_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111110111011101000100000001111111011101000100010000000000011111111111011101110100010000000111111101110100010001000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_11_S_1_out, I0 =>  C_11_S_1_L_0_out, I1 =>  C_11_S_1_L_1_out, I2 =>  C_11_S_1_L_2_out, I3 =>  C_11_S_1_L_3_out, I4 =>  C_11_S_1_L_4_out, I5 =>  C_11_S_1_L_5_out, I6 =>  C_11_S_1_L_6_out, I7 =>  C_11_S_1_L_7_out); 
C_11_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_11_S_2_out, I0 =>  C_11_S_2_L_0_out, I1 =>  C_11_S_2_L_1_out, I2 =>  C_11_S_2_L_2_out, I3 =>  C_11_S_2_L_3_out, I4 =>  C_11_S_2_L_4_out, I5 =>  C_11_S_2_L_5_out, I6 =>  C_11_S_2_L_6_out, I7 =>  C_11_S_2_L_7_out); 
C_11_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111111111011111110111010001111100011100000100000000000000011111111111111101111100011100000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_11_S_3_out, I0 =>  C_11_S_3_L_0_out, I1 =>  C_11_S_3_L_1_out, I2 =>  C_11_S_3_L_2_out, I3 =>  C_11_S_3_L_3_out, I4 =>  C_11_S_3_L_4_out, I5 =>  C_11_S_3_L_5_out, I6 =>  C_11_S_3_L_6_out, I7 =>  C_11_S_3_L_7_out); 
C_11_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111111111111011111110111010001111111010100000111111101110100011111000100000001110100010000000100000000000000011111111111111101111111011101000111111101110000011101000100000001111101010000000111010001000000010000000000000001000000000000000") port map( O =>C_11_S_4_out, I0 =>  C_11_S_4_L_0_out, I1 =>  C_11_S_4_L_1_out, I2 =>  C_11_S_4_L_2_out, I3 =>  C_11_S_4_L_3_out, I4 =>  C_11_S_4_L_4_out, I5 =>  C_11_S_4_L_5_out, I6 =>  C_11_S_4_L_6_out, I7 =>  C_11_S_4_L_7_out); 

C_11_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_11_out, I0 =>  C_11_S_0_out, I1 =>  C_11_S_1_out, I2 =>  C_11_S_2_out, I3 =>  C_11_S_3_out, I4 =>  C_11_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_12_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_12_S_0_out, I0 =>  C_12_S_0_L_0_out, I1 =>  C_12_S_0_L_1_out, I2 =>  C_12_S_0_L_2_out, I3 =>  C_12_S_0_L_3_out, I4 =>  C_12_S_0_L_4_out, I5 =>  C_12_S_0_L_5_out, I6 =>  C_12_S_0_L_6_out, I7 =>  C_12_S_0_L_7_out); 
C_12_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_12_S_1_out, I0 =>  C_12_S_1_L_0_out, I1 =>  C_12_S_1_L_1_out, I2 =>  C_12_S_1_L_2_out, I3 =>  C_12_S_1_L_3_out, I4 =>  C_12_S_1_L_4_out, I5 =>  C_12_S_1_L_5_out, I6 =>  C_12_S_1_L_6_out, I7 =>  C_12_S_1_L_7_out); 
C_12_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_12_S_2_out, I0 =>  C_12_S_2_L_0_out, I1 =>  C_12_S_2_L_1_out, I2 =>  C_12_S_2_L_2_out, I3 =>  C_12_S_2_L_3_out, I4 =>  C_12_S_2_L_4_out, I5 =>  C_12_S_2_L_5_out, I6 =>  C_12_S_2_L_6_out, I7 =>  C_12_S_2_L_7_out); 
C_12_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_12_S_3_out, I0 =>  C_12_S_3_L_0_out, I1 =>  C_12_S_3_L_1_out, I2 =>  C_12_S_3_L_2_out, I3 =>  C_12_S_3_L_3_out, I4 =>  C_12_S_3_L_4_out, I5 =>  C_12_S_3_L_5_out, I6 =>  C_12_S_3_L_6_out, I7 =>  C_12_S_3_L_7_out); 
C_12_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_12_S_4_out, I0 =>  C_12_S_4_L_0_out, I1 =>  C_12_S_4_L_1_out, I2 =>  C_12_S_4_L_2_out, I3 =>  C_12_S_4_L_3_out, I4 =>  C_12_S_4_L_4_out, I5 =>  C_12_S_4_L_5_out, I6 =>  C_12_S_4_L_6_out, I7 =>  C_12_S_4_L_7_out); 

C_12_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_12_out, I0 =>  C_12_S_0_out, I1 =>  C_12_S_1_out, I2 =>  C_12_S_2_out, I3 =>  C_12_S_3_out, I4 =>  C_12_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_13_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_13_S_0_out, I0 =>  C_13_S_0_L_0_out, I1 =>  C_13_S_0_L_1_out, I2 =>  C_13_S_0_L_2_out, I3 =>  C_13_S_0_L_3_out, I4 =>  C_13_S_0_L_4_out, I5 =>  C_13_S_0_L_5_out, I6 =>  C_13_S_0_L_6_out, I7 =>  C_13_S_0_L_7_out); 
C_13_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_13_S_1_out, I0 =>  C_13_S_1_L_0_out, I1 =>  C_13_S_1_L_1_out, I2 =>  C_13_S_1_L_2_out, I3 =>  C_13_S_1_L_3_out, I4 =>  C_13_S_1_L_4_out, I5 =>  C_13_S_1_L_5_out, I6 =>  C_13_S_1_L_6_out, I7 =>  C_13_S_1_L_7_out); 
C_13_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_13_S_2_out, I0 =>  C_13_S_2_L_0_out, I1 =>  C_13_S_2_L_1_out, I2 =>  C_13_S_2_L_2_out, I3 =>  C_13_S_2_L_3_out, I4 =>  C_13_S_2_L_4_out, I5 =>  C_13_S_2_L_5_out, I6 =>  C_13_S_2_L_6_out, I7 =>  C_13_S_2_L_7_out); 
C_13_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_13_S_3_out, I0 =>  C_13_S_3_L_0_out, I1 =>  C_13_S_3_L_1_out, I2 =>  C_13_S_3_L_2_out, I3 =>  C_13_S_3_L_3_out, I4 =>  C_13_S_3_L_4_out, I5 =>  C_13_S_3_L_5_out, I6 =>  C_13_S_3_L_6_out, I7 =>  C_13_S_3_L_7_out); 
C_13_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_13_S_4_out, I0 =>  C_13_S_4_L_0_out, I1 =>  C_13_S_4_L_1_out, I2 =>  C_13_S_4_L_2_out, I3 =>  C_13_S_4_L_3_out, I4 =>  C_13_S_4_L_4_out, I5 =>  C_13_S_4_L_5_out, I6 =>  C_13_S_4_L_6_out, I7 =>  C_13_S_4_L_7_out); 

C_13_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_13_out, I0 =>  C_13_S_0_out, I1 =>  C_13_S_1_out, I2 =>  C_13_S_2_out, I3 =>  C_13_S_3_out, I4 =>  C_13_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_14_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_14_S_0_out, I0 =>  C_14_S_0_L_0_out, I1 =>  C_14_S_0_L_1_out, I2 =>  C_14_S_0_L_2_out, I3 =>  C_14_S_0_L_3_out, I4 =>  C_14_S_0_L_4_out, I5 =>  C_14_S_0_L_5_out, I6 =>  C_14_S_0_L_6_out, I7 =>  C_14_S_0_L_7_out); 
C_14_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_14_S_1_out, I0 =>  C_14_S_1_L_0_out, I1 =>  C_14_S_1_L_1_out, I2 =>  C_14_S_1_L_2_out, I3 =>  C_14_S_1_L_3_out, I4 =>  C_14_S_1_L_4_out, I5 =>  C_14_S_1_L_5_out, I6 =>  C_14_S_1_L_6_out, I7 =>  C_14_S_1_L_7_out); 
C_14_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_14_S_2_out, I0 =>  C_14_S_2_L_0_out, I1 =>  C_14_S_2_L_1_out, I2 =>  C_14_S_2_L_2_out, I3 =>  C_14_S_2_L_3_out, I4 =>  C_14_S_2_L_4_out, I5 =>  C_14_S_2_L_5_out, I6 =>  C_14_S_2_L_6_out, I7 =>  C_14_S_2_L_7_out); 
C_14_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_14_S_3_out, I0 =>  C_14_S_3_L_0_out, I1 =>  C_14_S_3_L_1_out, I2 =>  C_14_S_3_L_2_out, I3 =>  C_14_S_3_L_3_out, I4 =>  C_14_S_3_L_4_out, I5 =>  C_14_S_3_L_5_out, I6 =>  C_14_S_3_L_6_out, I7 =>  C_14_S_3_L_7_out); 
C_14_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_14_S_4_out, I0 =>  C_14_S_4_L_0_out, I1 =>  C_14_S_4_L_1_out, I2 =>  C_14_S_4_L_2_out, I3 =>  C_14_S_4_L_3_out, I4 =>  C_14_S_4_L_4_out, I5 =>  C_14_S_4_L_5_out, I6 =>  C_14_S_4_L_6_out, I7 =>  C_14_S_4_L_7_out); 

C_14_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_14_out, I0 =>  C_14_S_0_out, I1 =>  C_14_S_1_out, I2 =>  C_14_S_2_out, I3 =>  C_14_S_3_out, I4 =>  C_14_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_15_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_15_S_0_out, I0 =>  C_15_S_0_L_0_out, I1 =>  C_15_S_0_L_1_out, I2 =>  C_15_S_0_L_2_out, I3 =>  C_15_S_0_L_3_out, I4 =>  C_15_S_0_L_4_out, I5 =>  C_15_S_0_L_5_out, I6 =>  C_15_S_0_L_6_out, I7 =>  C_15_S_0_L_7_out); 
C_15_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_15_S_1_out, I0 =>  C_15_S_1_L_0_out, I1 =>  C_15_S_1_L_1_out, I2 =>  C_15_S_1_L_2_out, I3 =>  C_15_S_1_L_3_out, I4 =>  C_15_S_1_L_4_out, I5 =>  C_15_S_1_L_5_out, I6 =>  C_15_S_1_L_6_out, I7 =>  C_15_S_1_L_7_out); 
C_15_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_15_S_2_out, I0 =>  C_15_S_2_L_0_out, I1 =>  C_15_S_2_L_1_out, I2 =>  C_15_S_2_L_2_out, I3 =>  C_15_S_2_L_3_out, I4 =>  C_15_S_2_L_4_out, I5 =>  C_15_S_2_L_5_out, I6 =>  C_15_S_2_L_6_out, I7 =>  C_15_S_2_L_7_out); 
C_15_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_15_S_3_out, I0 =>  C_15_S_3_L_0_out, I1 =>  C_15_S_3_L_1_out, I2 =>  C_15_S_3_L_2_out, I3 =>  C_15_S_3_L_3_out, I4 =>  C_15_S_3_L_4_out, I5 =>  C_15_S_3_L_5_out, I6 =>  C_15_S_3_L_6_out, I7 =>  C_15_S_3_L_7_out); 
C_15_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_15_S_4_out, I0 =>  C_15_S_4_L_0_out, I1 =>  C_15_S_4_L_1_out, I2 =>  C_15_S_4_L_2_out, I3 =>  C_15_S_4_L_3_out, I4 =>  C_15_S_4_L_4_out, I5 =>  C_15_S_4_L_5_out, I6 =>  C_15_S_4_L_6_out, I7 =>  C_15_S_4_L_7_out); 

C_15_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_15_out, I0 =>  C_15_S_0_out, I1 =>  C_15_S_1_out, I2 =>  C_15_S_2_out, I3 =>  C_15_S_3_out, I4 =>  C_15_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_16_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_16_S_0_out, I0 =>  C_16_S_0_L_0_out, I1 =>  C_16_S_0_L_1_out, I2 =>  C_16_S_0_L_2_out, I3 =>  C_16_S_0_L_3_out, I4 =>  C_16_S_0_L_4_out, I5 =>  C_16_S_0_L_5_out, I6 =>  C_16_S_0_L_6_out, I7 =>  C_16_S_0_L_7_out); 
C_16_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_16_S_1_out, I0 =>  C_16_S_1_L_0_out, I1 =>  C_16_S_1_L_1_out, I2 =>  C_16_S_1_L_2_out, I3 =>  C_16_S_1_L_3_out, I4 =>  C_16_S_1_L_4_out, I5 =>  C_16_S_1_L_5_out, I6 =>  C_16_S_1_L_6_out, I7 =>  C_16_S_1_L_7_out); 
C_16_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_16_S_2_out, I0 =>  C_16_S_2_L_0_out, I1 =>  C_16_S_2_L_1_out, I2 =>  C_16_S_2_L_2_out, I3 =>  C_16_S_2_L_3_out, I4 =>  C_16_S_2_L_4_out, I5 =>  C_16_S_2_L_5_out, I6 =>  C_16_S_2_L_6_out, I7 =>  C_16_S_2_L_7_out); 
C_16_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_16_S_3_out, I0 =>  C_16_S_3_L_0_out, I1 =>  C_16_S_3_L_1_out, I2 =>  C_16_S_3_L_2_out, I3 =>  C_16_S_3_L_3_out, I4 =>  C_16_S_3_L_4_out, I5 =>  C_16_S_3_L_5_out, I6 =>  C_16_S_3_L_6_out, I7 =>  C_16_S_3_L_7_out); 
C_16_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_16_S_4_out, I0 =>  C_16_S_4_L_0_out, I1 =>  C_16_S_4_L_1_out, I2 =>  C_16_S_4_L_2_out, I3 =>  C_16_S_4_L_3_out, I4 =>  C_16_S_4_L_4_out, I5 =>  C_16_S_4_L_5_out, I6 =>  C_16_S_4_L_6_out, I7 =>  C_16_S_4_L_7_out); 

C_16_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_16_out, I0 =>  C_16_S_0_out, I1 =>  C_16_S_1_out, I2 =>  C_16_S_2_out, I3 =>  C_16_S_3_out, I4 =>  C_16_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_17_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_17_S_0_out, I0 =>  C_17_S_0_L_0_out, I1 =>  C_17_S_0_L_1_out, I2 =>  C_17_S_0_L_2_out, I3 =>  C_17_S_0_L_3_out, I4 =>  C_17_S_0_L_4_out, I5 =>  C_17_S_0_L_5_out, I6 =>  C_17_S_0_L_6_out, I7 =>  C_17_S_0_L_7_out); 
C_17_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_17_S_1_out, I0 =>  C_17_S_1_L_0_out, I1 =>  C_17_S_1_L_1_out, I2 =>  C_17_S_1_L_2_out, I3 =>  C_17_S_1_L_3_out, I4 =>  C_17_S_1_L_4_out, I5 =>  C_17_S_1_L_5_out, I6 =>  C_17_S_1_L_6_out, I7 =>  C_17_S_1_L_7_out); 
C_17_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_17_S_2_out, I0 =>  C_17_S_2_L_0_out, I1 =>  C_17_S_2_L_1_out, I2 =>  C_17_S_2_L_2_out, I3 =>  C_17_S_2_L_3_out, I4 =>  C_17_S_2_L_4_out, I5 =>  C_17_S_2_L_5_out, I6 =>  C_17_S_2_L_6_out, I7 =>  C_17_S_2_L_7_out); 
C_17_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_17_S_3_out, I0 =>  C_17_S_3_L_0_out, I1 =>  C_17_S_3_L_1_out, I2 =>  C_17_S_3_L_2_out, I3 =>  C_17_S_3_L_3_out, I4 =>  C_17_S_3_L_4_out, I5 =>  C_17_S_3_L_5_out, I6 =>  C_17_S_3_L_6_out, I7 =>  C_17_S_3_L_7_out); 
C_17_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_17_S_4_out, I0 =>  C_17_S_4_L_0_out, I1 =>  C_17_S_4_L_1_out, I2 =>  C_17_S_4_L_2_out, I3 =>  C_17_S_4_L_3_out, I4 =>  C_17_S_4_L_4_out, I5 =>  C_17_S_4_L_5_out, I6 =>  C_17_S_4_L_6_out, I7 =>  C_17_S_4_L_7_out); 

C_17_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_17_out, I0 =>  C_17_S_0_out, I1 =>  C_17_S_1_out, I2 =>  C_17_S_2_out, I3 =>  C_17_S_3_out, I4 =>  C_17_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_18_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111010000000111111111111111011111110100000001111111010000000100000000000000011111111111111101111111010000000111111101000000010000000000000001111111010000000100000000000000010000000000000000000000000000000") port map( O =>C_18_S_0_out, I0 =>  C_18_S_0_L_0_out, I1 =>  C_18_S_0_L_1_out, I2 =>  C_18_S_0_L_2_out, I3 =>  C_18_S_0_L_3_out, I4 =>  C_18_S_0_L_4_out, I5 =>  C_18_S_0_L_5_out, I6 =>  C_18_S_0_L_6_out, I7 =>  C_18_S_0_L_7_out); 
C_18_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011100000111111111111111011111110111010001111111011101000111010000000000011111111111010001110100010000000111010001000000010000000000000001111100010000000100000000000000010000000000000000000000000000000") port map( O =>C_18_S_1_out, I0 =>  C_18_S_1_L_0_out, I1 =>  C_18_S_1_L_1_out, I2 =>  C_18_S_1_L_2_out, I3 =>  C_18_S_1_L_3_out, I4 =>  C_18_S_1_L_4_out, I5 =>  C_18_S_1_L_5_out, I6 =>  C_18_S_1_L_6_out, I7 =>  C_18_S_1_L_7_out); 
C_18_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_18_S_2_out, I0 =>  C_18_S_2_L_0_out, I1 =>  C_18_S_2_L_1_out, I2 =>  C_18_S_2_L_2_out, I3 =>  C_18_S_2_L_3_out, I4 =>  C_18_S_2_L_4_out, I5 =>  C_18_S_2_L_5_out, I6 =>  C_18_S_2_L_6_out, I7 =>  C_18_S_2_L_7_out); 
C_18_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111111111011111110111010001110100010000000100000000000000011111111111111101111111011101000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_18_S_3_out, I0 =>  C_18_S_3_L_0_out, I1 =>  C_18_S_3_L_1_out, I2 =>  C_18_S_3_L_2_out, I3 =>  C_18_S_3_L_3_out, I4 =>  C_18_S_3_L_4_out, I5 =>  C_18_S_3_L_5_out, I6 =>  C_18_S_3_L_6_out, I7 =>  C_18_S_3_L_7_out); 
C_18_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111101010000000111111111111111011111110101000001111111011101000101000000000000011111111111110101110100010000000111110101000000010000000000000001111111010100000100000000000000010000000000000000000000000000000") port map( O =>C_18_S_4_out, I0 =>  C_18_S_4_L_0_out, I1 =>  C_18_S_4_L_1_out, I2 =>  C_18_S_4_L_2_out, I3 =>  C_18_S_4_L_3_out, I4 =>  C_18_S_4_L_4_out, I5 =>  C_18_S_4_L_5_out, I6 =>  C_18_S_4_L_6_out, I7 =>  C_18_S_4_L_7_out); 

C_18_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_18_out, I0 =>  C_18_S_0_out, I1 =>  C_18_S_1_out, I2 =>  C_18_S_2_out, I3 =>  C_18_S_3_out, I4 =>  C_18_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_19_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_19_S_0_out, I0 =>  C_19_S_0_L_0_out, I1 =>  C_19_S_0_L_1_out, I2 =>  C_19_S_0_L_2_out, I3 =>  C_19_S_0_L_3_out, I4 =>  C_19_S_0_L_4_out, I5 =>  C_19_S_0_L_5_out, I6 =>  C_19_S_0_L_6_out, I7 =>  C_19_S_0_L_7_out); 
C_19_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_19_S_1_out, I0 =>  C_19_S_1_L_0_out, I1 =>  C_19_S_1_L_1_out, I2 =>  C_19_S_1_L_2_out, I3 =>  C_19_S_1_L_3_out, I4 =>  C_19_S_1_L_4_out, I5 =>  C_19_S_1_L_5_out, I6 =>  C_19_S_1_L_6_out, I7 =>  C_19_S_1_L_7_out); 
C_19_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_19_S_2_out, I0 =>  C_19_S_2_L_0_out, I1 =>  C_19_S_2_L_1_out, I2 =>  C_19_S_2_L_2_out, I3 =>  C_19_S_2_L_3_out, I4 =>  C_19_S_2_L_4_out, I5 =>  C_19_S_2_L_5_out, I6 =>  C_19_S_2_L_6_out, I7 =>  C_19_S_2_L_7_out); 
C_19_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_19_S_3_out, I0 =>  C_19_S_3_L_0_out, I1 =>  C_19_S_3_L_1_out, I2 =>  C_19_S_3_L_2_out, I3 =>  C_19_S_3_L_3_out, I4 =>  C_19_S_3_L_4_out, I5 =>  C_19_S_3_L_5_out, I6 =>  C_19_S_3_L_6_out, I7 =>  C_19_S_3_L_7_out); 
C_19_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_19_S_4_out, I0 =>  C_19_S_4_L_0_out, I1 =>  C_19_S_4_L_1_out, I2 =>  C_19_S_4_L_2_out, I3 =>  C_19_S_4_L_3_out, I4 =>  C_19_S_4_L_4_out, I5 =>  C_19_S_4_L_5_out, I6 =>  C_19_S_4_L_6_out, I7 =>  C_19_S_4_L_7_out); 

C_19_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_19_out, I0 =>  C_19_S_0_out, I1 =>  C_19_S_1_out, I2 =>  C_19_S_2_out, I3 =>  C_19_S_3_out, I4 =>  C_19_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_20_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_20_S_0_out, I0 =>  C_20_S_0_L_0_out, I1 =>  C_20_S_0_L_1_out, I2 =>  C_20_S_0_L_2_out, I3 =>  C_20_S_0_L_3_out, I4 =>  C_20_S_0_L_4_out, I5 =>  C_20_S_0_L_5_out, I6 =>  C_20_S_0_L_6_out, I7 =>  C_20_S_0_L_7_out); 
C_20_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_20_S_1_out, I0 =>  C_20_S_1_L_0_out, I1 =>  C_20_S_1_L_1_out, I2 =>  C_20_S_1_L_2_out, I3 =>  C_20_S_1_L_3_out, I4 =>  C_20_S_1_L_4_out, I5 =>  C_20_S_1_L_5_out, I6 =>  C_20_S_1_L_6_out, I7 =>  C_20_S_1_L_7_out); 
C_20_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_20_S_2_out, I0 =>  C_20_S_2_L_0_out, I1 =>  C_20_S_2_L_1_out, I2 =>  C_20_S_2_L_2_out, I3 =>  C_20_S_2_L_3_out, I4 =>  C_20_S_2_L_4_out, I5 =>  C_20_S_2_L_5_out, I6 =>  C_20_S_2_L_6_out, I7 =>  C_20_S_2_L_7_out); 
C_20_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_20_S_3_out, I0 =>  C_20_S_3_L_0_out, I1 =>  C_20_S_3_L_1_out, I2 =>  C_20_S_3_L_2_out, I3 =>  C_20_S_3_L_3_out, I4 =>  C_20_S_3_L_4_out, I5 =>  C_20_S_3_L_5_out, I6 =>  C_20_S_3_L_6_out, I7 =>  C_20_S_3_L_7_out); 
C_20_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_20_S_4_out, I0 =>  C_20_S_4_L_0_out, I1 =>  C_20_S_4_L_1_out, I2 =>  C_20_S_4_L_2_out, I3 =>  C_20_S_4_L_3_out, I4 =>  C_20_S_4_L_4_out, I5 =>  C_20_S_4_L_5_out, I6 =>  C_20_S_4_L_6_out, I7 =>  C_20_S_4_L_7_out); 

C_20_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_20_out, I0 =>  C_20_S_0_out, I1 =>  C_20_S_1_out, I2 =>  C_20_S_2_out, I3 =>  C_20_S_3_out, I4 =>  C_20_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_21_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111010000000111111111111111011111110100000001111111010000000100000000000000011111111111111101111111010000000111111101000000010000000000000001111111010000000100000000000000010000000000000000000000000000000") port map( O =>C_21_S_0_out, I0 =>  C_21_S_0_L_0_out, I1 =>  C_21_S_0_L_1_out, I2 =>  C_21_S_0_L_2_out, I3 =>  C_21_S_0_L_3_out, I4 =>  C_21_S_0_L_4_out, I5 =>  C_21_S_0_L_5_out, I6 =>  C_21_S_0_L_6_out, I7 =>  C_21_S_0_L_7_out); 
C_21_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011100000111111111111111011111110111010001111111011101000111010000000000011111111111010001110100010000000111010001000000010000000000000001111100010000000100000000000000010000000000000000000000000000000") port map( O =>C_21_S_1_out, I0 =>  C_21_S_1_L_0_out, I1 =>  C_21_S_1_L_1_out, I2 =>  C_21_S_1_L_2_out, I3 =>  C_21_S_1_L_3_out, I4 =>  C_21_S_1_L_4_out, I5 =>  C_21_S_1_L_5_out, I6 =>  C_21_S_1_L_6_out, I7 =>  C_21_S_1_L_7_out); 
C_21_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_21_S_2_out, I0 =>  C_21_S_2_L_0_out, I1 =>  C_21_S_2_L_1_out, I2 =>  C_21_S_2_L_2_out, I3 =>  C_21_S_2_L_3_out, I4 =>  C_21_S_2_L_4_out, I5 =>  C_21_S_2_L_5_out, I6 =>  C_21_S_2_L_6_out, I7 =>  C_21_S_2_L_7_out); 
C_21_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111111111011111110111010001110100010000000100000000000000011111111111111101111111011101000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_21_S_3_out, I0 =>  C_21_S_3_L_0_out, I1 =>  C_21_S_3_L_1_out, I2 =>  C_21_S_3_L_2_out, I3 =>  C_21_S_3_L_3_out, I4 =>  C_21_S_3_L_4_out, I5 =>  C_21_S_3_L_5_out, I6 =>  C_21_S_3_L_6_out, I7 =>  C_21_S_3_L_7_out); 
C_21_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111101010000000111111111111111011111110101000001111111011101000101000000000000011111111111110101110100010000000111110101000000010000000000000001111111010100000100000000000000010000000000000000000000000000000") port map( O =>C_21_S_4_out, I0 =>  C_21_S_4_L_0_out, I1 =>  C_21_S_4_L_1_out, I2 =>  C_21_S_4_L_2_out, I3 =>  C_21_S_4_L_3_out, I4 =>  C_21_S_4_L_4_out, I5 =>  C_21_S_4_L_5_out, I6 =>  C_21_S_4_L_6_out, I7 =>  C_21_S_4_L_7_out); 

C_21_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_21_out, I0 =>  C_21_S_0_out, I1 =>  C_21_S_1_out, I2 =>  C_21_S_2_out, I3 =>  C_21_S_3_out, I4 =>  C_21_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_22_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_22_S_0_out, I0 =>  C_22_S_0_L_0_out, I1 =>  C_22_S_0_L_1_out, I2 =>  C_22_S_0_L_2_out, I3 =>  C_22_S_0_L_3_out, I4 =>  C_22_S_0_L_4_out, I5 =>  C_22_S_0_L_5_out, I6 =>  C_22_S_0_L_6_out, I7 =>  C_22_S_0_L_7_out); 
C_22_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_22_S_1_out, I0 =>  C_22_S_1_L_0_out, I1 =>  C_22_S_1_L_1_out, I2 =>  C_22_S_1_L_2_out, I3 =>  C_22_S_1_L_3_out, I4 =>  C_22_S_1_L_4_out, I5 =>  C_22_S_1_L_5_out, I6 =>  C_22_S_1_L_6_out, I7 =>  C_22_S_1_L_7_out); 
C_22_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_22_S_2_out, I0 =>  C_22_S_2_L_0_out, I1 =>  C_22_S_2_L_1_out, I2 =>  C_22_S_2_L_2_out, I3 =>  C_22_S_2_L_3_out, I4 =>  C_22_S_2_L_4_out, I5 =>  C_22_S_2_L_5_out, I6 =>  C_22_S_2_L_6_out, I7 =>  C_22_S_2_L_7_out); 
C_22_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_22_S_3_out, I0 =>  C_22_S_3_L_0_out, I1 =>  C_22_S_3_L_1_out, I2 =>  C_22_S_3_L_2_out, I3 =>  C_22_S_3_L_3_out, I4 =>  C_22_S_3_L_4_out, I5 =>  C_22_S_3_L_5_out, I6 =>  C_22_S_3_L_6_out, I7 =>  C_22_S_3_L_7_out); 
C_22_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_22_S_4_out, I0 =>  C_22_S_4_L_0_out, I1 =>  C_22_S_4_L_1_out, I2 =>  C_22_S_4_L_2_out, I3 =>  C_22_S_4_L_3_out, I4 =>  C_22_S_4_L_4_out, I5 =>  C_22_S_4_L_5_out, I6 =>  C_22_S_4_L_6_out, I7 =>  C_22_S_4_L_7_out); 

C_22_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_22_out, I0 =>  C_22_S_0_out, I1 =>  C_22_S_1_out, I2 =>  C_22_S_2_out, I3 =>  C_22_S_3_out, I4 =>  C_22_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_23_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_23_S_0_out, I0 =>  C_23_S_0_L_0_out, I1 =>  C_23_S_0_L_1_out, I2 =>  C_23_S_0_L_2_out, I3 =>  C_23_S_0_L_3_out, I4 =>  C_23_S_0_L_4_out, I5 =>  C_23_S_0_L_5_out, I6 =>  C_23_S_0_L_6_out, I7 =>  C_23_S_0_L_7_out); 
C_23_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_23_S_1_out, I0 =>  C_23_S_1_L_0_out, I1 =>  C_23_S_1_L_1_out, I2 =>  C_23_S_1_L_2_out, I3 =>  C_23_S_1_L_3_out, I4 =>  C_23_S_1_L_4_out, I5 =>  C_23_S_1_L_5_out, I6 =>  C_23_S_1_L_6_out, I7 =>  C_23_S_1_L_7_out); 
C_23_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_23_S_2_out, I0 =>  C_23_S_2_L_0_out, I1 =>  C_23_S_2_L_1_out, I2 =>  C_23_S_2_L_2_out, I3 =>  C_23_S_2_L_3_out, I4 =>  C_23_S_2_L_4_out, I5 =>  C_23_S_2_L_5_out, I6 =>  C_23_S_2_L_6_out, I7 =>  C_23_S_2_L_7_out); 
C_23_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_23_S_3_out, I0 =>  C_23_S_3_L_0_out, I1 =>  C_23_S_3_L_1_out, I2 =>  C_23_S_3_L_2_out, I3 =>  C_23_S_3_L_3_out, I4 =>  C_23_S_3_L_4_out, I5 =>  C_23_S_3_L_5_out, I6 =>  C_23_S_3_L_6_out, I7 =>  C_23_S_3_L_7_out); 
C_23_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111101011111111111110101111101010100000111111111111101011111010101000001111101010100000101000000000000011111111111110101111101010100000111110101010000010100000000000001111101010100000101000000000000010100000000000000000000000000000") port map( O =>C_23_S_4_out, I0 =>  C_23_S_4_L_0_out, I1 =>  C_23_S_4_L_1_out, I2 =>  C_23_S_4_L_2_out, I3 =>  C_23_S_4_L_3_out, I4 =>  C_23_S_4_L_4_out, I5 =>  C_23_S_4_L_5_out, I6 =>  C_23_S_4_L_6_out, I7 =>  C_23_S_4_L_7_out); 

C_23_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_23_out, I0 =>  C_23_S_0_out, I1 =>  C_23_S_1_out, I2 =>  C_23_S_2_out, I3 =>  C_23_S_3_out, I4 =>  C_23_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_24_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101000111011101110101011101010101010101110101010101010101010101010100011101010101010101010101010101000101010101010100010101000100010001110101010101010101010101010100010101010101010001010100010000000") port map( O =>C_24_S_0_out, I0 =>  C_24_S_0_L_0_out, I1 =>  C_24_S_0_L_1_out, I2 =>  C_24_S_0_L_2_out, I3 =>  C_24_S_0_L_3_out, I4 =>  C_24_S_0_L_4_out, I5 =>  C_24_S_0_L_5_out, I6 =>  C_24_S_0_L_6_out, I7 =>  C_24_S_0_L_7_out); 
C_24_S_1_inst : LUT8 generic map(INIT => "1111111111111100111111101110100011111110111010001111100011100000111111101110100011111000111000001111110011100000111010001000000011111110111010001111100011000000111110001110000011101000100000001111100011100000111010001000000011101000100000001100000000000000") port map( O =>C_24_S_1_out, I0 =>  C_24_S_1_L_0_out, I1 =>  C_24_S_1_L_1_out, I2 =>  C_24_S_1_L_2_out, I3 =>  C_24_S_1_L_3_out, I4 =>  C_24_S_1_L_4_out, I5 =>  C_24_S_1_L_5_out, I6 =>  C_24_S_1_L_6_out, I7 =>  C_24_S_1_L_7_out); 
C_24_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111110101011111111111111101110111010101000111111101110100011101000100000001110101010000000100000000000000011111111111111101111111010101000111111101110100011101000100000001110101010001000100000000000000010101000000000000000000000000000") port map( O =>C_24_S_2_out, I0 =>  C_24_S_2_L_0_out, I1 =>  C_24_S_2_L_1_out, I2 =>  C_24_S_2_L_2_out, I3 =>  C_24_S_2_L_3_out, I4 =>  C_24_S_2_L_4_out, I5 =>  C_24_S_2_L_5_out, I6 =>  C_24_S_2_L_6_out, I7 =>  C_24_S_2_L_7_out); 
C_24_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110111010000000111111101110100011101000100000001110100010000000100010000000000011111111111011101111111011101000111111101110100011101000100000001111111010001000111010001000000011101000100000001000000000000000") port map( O =>C_24_S_3_out, I0 =>  C_24_S_3_L_0_out, I1 =>  C_24_S_3_L_1_out, I2 =>  C_24_S_3_L_2_out, I3 =>  C_24_S_3_L_3_out, I4 =>  C_24_S_3_L_4_out, I5 =>  C_24_S_3_L_5_out, I6 =>  C_24_S_3_L_6_out, I7 =>  C_24_S_3_L_7_out); 
C_24_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101111110011111111111111001111110011101000111111101111110011111100110000001111110011101000111010001000000011111110111010001110100011000000111111001100000011000000100000001110100011000000110000000000000011000000100000001000000000000000") port map( O =>C_24_S_4_out, I0 =>  C_24_S_4_L_0_out, I1 =>  C_24_S_4_L_1_out, I2 =>  C_24_S_4_L_2_out, I3 =>  C_24_S_4_L_3_out, I4 =>  C_24_S_4_L_4_out, I5 =>  C_24_S_4_L_5_out, I6 =>  C_24_S_4_L_6_out, I7 =>  C_24_S_4_L_7_out); 

C_24_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_24_out, I0 =>  C_24_S_0_out, I1 =>  C_24_S_1_out, I2 =>  C_24_S_2_out, I3 =>  C_24_S_3_out, I4 =>  C_24_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_25_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111110100010001110111010000000100000000000000011111111111111101111111010001000111011101000000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_25_S_0_out, I0 =>  C_25_S_0_L_0_out, I1 =>  C_25_S_0_L_1_out, I2 =>  C_25_S_0_L_2_out, I3 =>  C_25_S_0_L_3_out, I4 =>  C_25_S_0_L_4_out, I5 =>  C_25_S_0_L_5_out, I6 =>  C_25_S_0_L_6_out, I7 =>  C_25_S_0_L_7_out); 
C_25_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_25_S_1_out, I0 =>  C_25_S_1_L_0_out, I1 =>  C_25_S_1_L_1_out, I2 =>  C_25_S_1_L_2_out, I3 =>  C_25_S_1_L_3_out, I4 =>  C_25_S_1_L_4_out, I5 =>  C_25_S_1_L_5_out, I6 =>  C_25_S_1_L_6_out, I7 =>  C_25_S_1_L_7_out); 
C_25_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111111111010001110100010000000111111101110100011101000100000001111111011101000111010000000000011111111111010001110100010000000111111101110100011101000100000001111111011101000111010000000000011101000100000001000000000000000") port map( O =>C_25_S_2_out, I0 =>  C_25_S_2_L_0_out, I1 =>  C_25_S_2_L_1_out, I2 =>  C_25_S_2_L_2_out, I3 =>  C_25_S_2_L_3_out, I4 =>  C_25_S_2_L_4_out, I5 =>  C_25_S_2_L_5_out, I6 =>  C_25_S_2_L_6_out, I7 =>  C_25_S_2_L_7_out); 
C_25_S_3_inst : LUT8 generic map(INIT => "1111111111111010111111101110100011111110111010001111100010100000111111101110100011111000101000001111111011101000111010001000000011111110111010001110100010000000111110101110000011101000100000001111101011100000111010001000000011101000100000001010000000000000") port map( O =>C_25_S_3_out, I0 =>  C_25_S_3_L_0_out, I1 =>  C_25_S_3_L_1_out, I2 =>  C_25_S_3_L_2_out, I3 =>  C_25_S_3_L_3_out, I4 =>  C_25_S_3_L_4_out, I5 =>  C_25_S_3_L_5_out, I6 =>  C_25_S_3_L_6_out, I7 =>  C_25_S_3_L_7_out); 
C_25_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111101011111110111010001110100010000000111010000000000011111111111010001111111011101000111010001000000010100000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_25_S_4_out, I0 =>  C_25_S_4_L_0_out, I1 =>  C_25_S_4_L_1_out, I2 =>  C_25_S_4_L_2_out, I3 =>  C_25_S_4_L_3_out, I4 =>  C_25_S_4_L_4_out, I5 =>  C_25_S_4_L_5_out, I6 =>  C_25_S_4_L_6_out, I7 =>  C_25_S_4_L_7_out); 

C_25_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_25_out, I0 =>  C_25_S_0_out, I1 =>  C_25_S_1_out, I2 =>  C_25_S_2_out, I3 =>  C_25_S_3_out, I4 =>  C_25_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_26_S_0_inst : LUT8 generic map(INIT => "1111111011111110111110101110100011111010111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001010000011101000101000001000000010000000") port map( O =>C_26_S_0_out, I0 =>  C_26_S_0_L_0_out, I1 =>  C_26_S_0_L_1_out, I2 =>  C_26_S_0_L_2_out, I3 =>  C_26_S_0_L_3_out, I4 =>  C_26_S_0_L_4_out, I5 =>  C_26_S_0_L_5_out, I6 =>  C_26_S_0_L_6_out, I7 =>  C_26_S_0_L_7_out); 
C_26_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011101110111011101110111010101000111011101110100011101010100010001110100010001000100010001000000011111110111011101110111011101000111011101010100011101000100010001110101010001000100010001000100010001000100000001000000000000000") port map( O =>C_26_S_1_out, I0 =>  C_26_S_1_L_0_out, I1 =>  C_26_S_1_L_1_out, I2 =>  C_26_S_1_L_2_out, I3 =>  C_26_S_1_L_3_out, I4 =>  C_26_S_1_L_4_out, I5 =>  C_26_S_1_L_5_out, I6 =>  C_26_S_1_L_6_out, I7 =>  C_26_S_1_L_7_out); 
C_26_S_2_inst : LUT8 generic map(INIT => "1111111011111110111111101110101011111110111010101110111011101000111011101110100011101000101010001110101011101000111010001000000011111110111010001110100010101000111010101110100011101000100010001110100010001000101010001000000010101000100000001000000010000000") port map( O =>C_26_S_2_out, I0 =>  C_26_S_2_L_0_out, I1 =>  C_26_S_2_L_1_out, I2 =>  C_26_S_2_L_2_out, I3 =>  C_26_S_2_L_3_out, I4 =>  C_26_S_2_L_4_out, I5 =>  C_26_S_2_L_5_out, I6 =>  C_26_S_2_L_6_out, I7 =>  C_26_S_2_L_7_out); 
C_26_S_3_inst : LUT8 generic map(INIT => "1111111011101110111111101110101011101110111010101110101011101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110100010101000101010001000100010101000100000001000100010000000") port map( O =>C_26_S_3_out, I0 =>  C_26_S_3_L_0_out, I1 =>  C_26_S_3_L_1_out, I2 =>  C_26_S_3_L_2_out, I3 =>  C_26_S_3_L_3_out, I4 =>  C_26_S_3_L_4_out, I5 =>  C_26_S_3_L_5_out, I6 =>  C_26_S_3_L_6_out, I7 =>  C_26_S_3_L_7_out); 
C_26_S_4_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011111110111011101110111011101000111011101110100011101000101010001110101010101000111010001000100011101110111010001110101010101000111010101110100011101000100010001110100010001000100010001000000010101000100010001000100010000000") port map( O =>C_26_S_4_out, I0 =>  C_26_S_4_L_0_out, I1 =>  C_26_S_4_L_1_out, I2 =>  C_26_S_4_L_2_out, I3 =>  C_26_S_4_L_3_out, I4 =>  C_26_S_4_L_4_out, I5 =>  C_26_S_4_L_5_out, I6 =>  C_26_S_4_L_6_out, I7 =>  C_26_S_4_L_7_out); 

C_26_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_26_out, I0 =>  C_26_S_0_out, I1 =>  C_26_S_1_out, I2 =>  C_26_S_2_out, I3 =>  C_26_S_3_out, I4 =>  C_26_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_27_S_0_inst : LUT8 generic map(INIT => "1111111011101010111110101010101011101010101010101110101010101000111110101110101011101010101010001110101010101000101010101010000011111010101010101110101010101000111010101010100010101000101000001110101010101000101010101010100010101010101000001010100010000000") port map( O =>C_27_S_0_out, I0 =>  C_27_S_0_L_0_out, I1 =>  C_27_S_0_L_1_out, I2 =>  C_27_S_0_L_2_out, I3 =>  C_27_S_0_L_3_out, I4 =>  C_27_S_0_L_4_out, I5 =>  C_27_S_0_L_5_out, I6 =>  C_27_S_0_L_6_out, I7 =>  C_27_S_0_L_7_out); 
C_27_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110111010001000111111101110100011101110100010001110111010001000111010001000000011111110111010001110111010001000111011101000100011101000100000001110111010001000111010001000000011101000100000001000000000000000") port map( O =>C_27_S_1_out, I0 =>  C_27_S_1_L_0_out, I1 =>  C_27_S_1_L_1_out, I2 =>  C_27_S_1_L_2_out, I3 =>  C_27_S_1_L_3_out, I4 =>  C_27_S_1_L_4_out, I5 =>  C_27_S_1_L_5_out, I6 =>  C_27_S_1_L_6_out, I7 =>  C_27_S_1_L_7_out); 
C_27_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111101110101011111110111010101110101010101000111111101110101011101010101010001110101010101000100000000000000011111111111111101110101010101000111010101010100010101000100000001110101010101000101010001000000010101000100000000000000000000000") port map( O =>C_27_S_2_out, I0 =>  C_27_S_2_L_0_out, I1 =>  C_27_S_2_L_1_out, I2 =>  C_27_S_2_L_2_out, I3 =>  C_27_S_2_L_3_out, I4 =>  C_27_S_2_L_4_out, I5 =>  C_27_S_2_L_5_out, I6 =>  C_27_S_2_L_6_out, I7 =>  C_27_S_2_L_7_out); 
C_27_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111111110101011111110111010001111111011101000111111101110100011111110101010001110100010000000111010001000000011111110111010001111111011101000111010101000000011101000100000001110100010000000111010001000000010101000000000001000000000000000") port map( O =>C_27_S_3_out, I0 =>  C_27_S_3_L_0_out, I1 =>  C_27_S_3_L_1_out, I2 =>  C_27_S_3_L_2_out, I3 =>  C_27_S_3_L_3_out, I4 =>  C_27_S_3_L_4_out, I5 =>  C_27_S_3_L_5_out, I6 =>  C_27_S_3_L_6_out, I7 =>  C_27_S_3_L_7_out); 
C_27_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110110011111110111011001110110011001000111111101110110011101000110010001110100011001000100010001000000011111110111011101110110011101000111011001110100011001000100000001110110011001000110010001000000011001000100000001000000000000000") port map( O =>C_27_S_4_out, I0 =>  C_27_S_4_L_0_out, I1 =>  C_27_S_4_L_1_out, I2 =>  C_27_S_4_L_2_out, I3 =>  C_27_S_4_L_3_out, I4 =>  C_27_S_4_L_4_out, I5 =>  C_27_S_4_L_5_out, I6 =>  C_27_S_4_L_6_out, I7 =>  C_27_S_4_L_7_out); 

C_27_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_27_out, I0 =>  C_27_S_0_out, I1 =>  C_27_S_1_out, I2 =>  C_27_S_2_out, I3 =>  C_27_S_3_out, I4 =>  C_27_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_28_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101110101010101000111010101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000101010001110101010101000101010101010100010101010101010001010100010000000") port map( O =>C_28_S_0_out, I0 =>  C_28_S_0_L_0_out, I1 =>  C_28_S_0_L_1_out, I2 =>  C_28_S_0_L_2_out, I3 =>  C_28_S_0_L_3_out, I4 =>  C_28_S_0_L_4_out, I5 =>  C_28_S_0_L_5_out, I6 =>  C_28_S_0_L_6_out, I7 =>  C_28_S_0_L_7_out); 
C_28_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111111010101011111111111010101110101010000000111111111110101011101110100000001111111010000000101010000000000011111111111010101111111010000000111111101000100010101000000000001111111010101000101010000000000010101010000000001000000000000000") port map( O =>C_28_S_1_out, I0 =>  C_28_S_1_L_0_out, I1 =>  C_28_S_1_L_1_out, I2 =>  C_28_S_1_L_2_out, I3 =>  C_28_S_1_L_3_out, I4 =>  C_28_S_1_L_4_out, I5 =>  C_28_S_1_L_5_out, I6 =>  C_28_S_1_L_6_out, I7 =>  C_28_S_1_L_7_out); 
C_28_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101110101010001000111111111111111011101110111010001110111011101000100010001000000011111110111011101110100010001000111010001000100010000000000000001110111010101000100000000000000010000000000000000000000000000000") port map( O =>C_28_S_2_out, I0 =>  C_28_S_2_L_0_out, I1 =>  C_28_S_2_L_1_out, I2 =>  C_28_S_2_L_2_out, I3 =>  C_28_S_2_L_3_out, I4 =>  C_28_S_2_L_4_out, I5 =>  C_28_S_2_L_5_out, I6 =>  C_28_S_2_L_6_out, I7 =>  C_28_S_2_L_7_out); 
C_28_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101111111011111110111010001110100011100000111111101111111011111110111010001110100011100000100000001000000011111110111111101111100011101000111010001000000010000000100000001111100011101000111010001000000010000000100000001000000000000000") port map( O =>C_28_S_3_out, I0 =>  C_28_S_3_L_0_out, I1 =>  C_28_S_3_L_1_out, I2 =>  C_28_S_3_L_2_out, I3 =>  C_28_S_3_L_3_out, I4 =>  C_28_S_3_L_4_out, I5 =>  C_28_S_3_L_5_out, I6 =>  C_28_S_3_L_6_out, I7 =>  C_28_S_3_L_7_out); 
C_28_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101011101000111111101110100011101000100010001110100010101000101010001000000011111110111010101110101011101000111011101110100011101000100000001110100010101000101010001000000010101000100000001000000000000000") port map( O =>C_28_S_4_out, I0 =>  C_28_S_4_L_0_out, I1 =>  C_28_S_4_L_1_out, I2 =>  C_28_S_4_L_2_out, I3 =>  C_28_S_4_L_3_out, I4 =>  C_28_S_4_L_4_out, I5 =>  C_28_S_4_L_5_out, I6 =>  C_28_S_4_L_6_out, I7 =>  C_28_S_4_L_7_out); 

C_28_inst : LUT8 generic map(INIT => "1111100011101000111010001110000011111000111010001110100011100000111110001110100011101000111000001111100011101000111010001110000011111000111010001110100011100000111110001110100011101000111000001111100011101000111010001110000011111000111010001110100011100000") port map( O =>C_28_out, I0 =>  C_28_S_0_out, I1 =>  C_28_S_1_out, I2 =>  C_28_S_2_out, I3 =>  C_28_S_3_out, I4 =>  C_28_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_29_S_0_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010101110100010001000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110111011101000101010001000100011101000100010001000100010000000") port map( O =>C_29_S_0_out, I0 =>  C_29_S_0_L_0_out, I1 =>  C_29_S_0_L_1_out, I2 =>  C_29_S_0_L_2_out, I3 =>  C_29_S_0_L_3_out, I4 =>  C_29_S_0_L_4_out, I5 =>  C_29_S_0_L_5_out, I6 =>  C_29_S_0_L_6_out, I7 =>  C_29_S_0_L_7_out); 
C_29_S_1_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_29_S_1_out, I0 =>  C_29_S_1_L_0_out, I1 =>  C_29_S_1_L_1_out, I2 =>  C_29_S_1_L_2_out, I3 =>  C_29_S_1_L_3_out, I4 =>  C_29_S_1_L_4_out, I5 =>  C_29_S_1_L_5_out, I6 =>  C_29_S_1_L_6_out, I7 =>  C_29_S_1_L_7_out); 
C_29_S_2_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111111101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100000001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_29_S_2_out, I0 =>  C_29_S_2_L_0_out, I1 =>  C_29_S_2_L_1_out, I2 =>  C_29_S_2_L_2_out, I3 =>  C_29_S_2_L_3_out, I4 =>  C_29_S_2_L_4_out, I5 =>  C_29_S_2_L_5_out, I6 =>  C_29_S_2_L_6_out, I7 =>  C_29_S_2_L_7_out); 
C_29_S_3_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010101110100010001000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110111011101000101010001000100011101000100010001000100010000000") port map( O =>C_29_S_3_out, I0 =>  C_29_S_3_L_0_out, I1 =>  C_29_S_3_L_1_out, I2 =>  C_29_S_3_L_2_out, I3 =>  C_29_S_3_L_3_out, I4 =>  C_29_S_3_L_4_out, I5 =>  C_29_S_3_L_5_out, I6 =>  C_29_S_3_L_6_out, I7 =>  C_29_S_3_L_7_out); 
C_29_S_4_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_29_S_4_out, I0 =>  C_29_S_4_L_0_out, I1 =>  C_29_S_4_L_1_out, I2 =>  C_29_S_4_L_2_out, I3 =>  C_29_S_4_L_3_out, I4 =>  C_29_S_4_L_4_out, I5 =>  C_29_S_4_L_5_out, I6 =>  C_29_S_4_L_6_out, I7 =>  C_29_S_4_L_7_out); 

C_29_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_29_out, I0 =>  C_29_S_0_out, I1 =>  C_29_S_1_out, I2 =>  C_29_S_2_out, I3 =>  C_29_S_3_out, I4 =>  C_29_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_30_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101000111010101110101011101010101010001110101010101010101010101010100011101010101010101010101010101000111010101010100010101000101010001110101010101010101010101010100010101010101010001010100010000000") port map( O =>C_30_S_0_out, I0 =>  C_30_S_0_L_0_out, I1 =>  C_30_S_0_L_1_out, I2 =>  C_30_S_0_L_2_out, I3 =>  C_30_S_0_L_3_out, I4 =>  C_30_S_0_L_4_out, I5 =>  C_30_S_0_L_5_out, I6 =>  C_30_S_0_L_6_out, I7 =>  C_30_S_0_L_7_out); 
C_30_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011101110101010001110111010001000100010000000000011111111111011101110111010001000111010101000100010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_30_S_1_out, I0 =>  C_30_S_1_L_0_out, I1 =>  C_30_S_1_L_1_out, I2 =>  C_30_S_1_L_2_out, I3 =>  C_30_S_1_L_3_out, I4 =>  C_30_S_1_L_4_out, I5 =>  C_30_S_1_L_5_out, I6 =>  C_30_S_1_L_6_out, I7 =>  C_30_S_1_L_7_out); 
C_30_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110111010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010001000101010001000000010101000100000001000000000000000") port map( O =>C_30_S_2_out, I0 =>  C_30_S_2_L_0_out, I1 =>  C_30_S_2_L_1_out, I2 =>  C_30_S_2_L_2_out, I3 =>  C_30_S_2_L_3_out, I4 =>  C_30_S_2_L_4_out, I5 =>  C_30_S_2_L_5_out, I6 =>  C_30_S_2_L_6_out, I7 =>  C_30_S_2_L_7_out); 
C_30_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111111111110011111110111010001111110011000000111111111111110011111110111010001111110011000000111010001000000011111110111010001111110011000000111010001000000011000000000000001111110011000000111010001000000011000000000000001000000000000000") port map( O =>C_30_S_3_out, I0 =>  C_30_S_3_L_0_out, I1 =>  C_30_S_3_L_1_out, I2 =>  C_30_S_3_L_2_out, I3 =>  C_30_S_3_L_3_out, I4 =>  C_30_S_3_L_4_out, I5 =>  C_30_S_3_L_5_out, I6 =>  C_30_S_3_L_6_out, I7 =>  C_30_S_3_L_7_out); 
C_30_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111101110111011111110111011101110100010001000111111101110111011101110111010001110111011101000100010001000000011111110111011101110100010001000111010001000100010001000100000001110111011101000100010001000000010001000100000000000000000000000") port map( O =>C_30_S_4_out, I0 =>  C_30_S_4_L_0_out, I1 =>  C_30_S_4_L_1_out, I2 =>  C_30_S_4_L_2_out, I3 =>  C_30_S_4_L_3_out, I4 =>  C_30_S_4_L_4_out, I5 =>  C_30_S_4_L_5_out, I6 =>  C_30_S_4_L_6_out, I7 =>  C_30_S_4_L_7_out); 

C_30_inst : LUT8 generic map(INIT => "1110101011101000111010001010100011101010111010001110100010101000111010101110100011101000101010001110101011101000111010001010100011101010111010001110100010101000111010101110100011101000101010001110101011101000111010001010100011101010111010001110100010101000") port map( O =>C_30_out, I0 =>  C_30_S_0_out, I1 =>  C_30_S_1_out, I2 =>  C_30_S_2_out, I3 =>  C_30_S_3_out, I4 =>  C_30_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_31_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101010100011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100011101010101010001010100010000000") port map( O =>C_31_S_0_out, I0 =>  C_31_S_0_L_0_out, I1 =>  C_31_S_0_L_1_out, I2 =>  C_31_S_0_L_2_out, I3 =>  C_31_S_0_L_3_out, I4 =>  C_31_S_0_L_4_out, I5 =>  C_31_S_0_L_5_out, I6 =>  C_31_S_0_L_6_out, I7 =>  C_31_S_0_L_7_out); 
C_31_S_1_inst : LUT8 generic map(INIT => "1111111011101010111111101110101011111110111010101110101010101000111110101110101011101010101010001110101010101000101010101010000011111010101010101110101010101000111010101010100010101000101000001110101010101000101010001000000010101000100000001010100010000000") port map( O =>C_31_S_1_out, I0 =>  C_31_S_1_L_0_out, I1 =>  C_31_S_1_L_1_out, I2 =>  C_31_S_1_L_2_out, I3 =>  C_31_S_1_L_3_out, I4 =>  C_31_S_1_L_4_out, I5 =>  C_31_S_1_L_5_out, I6 =>  C_31_S_1_L_6_out, I7 =>  C_31_S_1_L_7_out); 
C_31_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111101111110011111110111110001111100011100000111111101111110011111000111000001111100011100000111000001000000011111110111110001111100011100000111110001110000011000000100000001111100011100000111000001000000011000000100000000000000000000000") port map( O =>C_31_S_2_out, I0 =>  C_31_S_2_L_0_out, I1 =>  C_31_S_2_L_1_out, I2 =>  C_31_S_2_L_2_out, I3 =>  C_31_S_2_L_3_out, I4 =>  C_31_S_2_L_4_out, I5 =>  C_31_S_2_L_5_out, I6 =>  C_31_S_2_L_6_out, I7 =>  C_31_S_2_L_7_out); 
C_31_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111101111111011111110111111001111100011101000111111101111100011101000111000001110100010000000100000001000000011111110111111101111111011101000111110001110100011100000100000001110100011100000110000001000000010000000100000000000000000000000") port map( O =>C_31_S_3_out, I0 =>  C_31_S_3_L_0_out, I1 =>  C_31_S_3_L_1_out, I2 =>  C_31_S_3_L_2_out, I3 =>  C_31_S_3_L_3_out, I4 =>  C_31_S_3_L_4_out, I5 =>  C_31_S_3_L_5_out, I6 =>  C_31_S_3_L_6_out, I7 =>  C_31_S_3_L_7_out); 
C_31_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111101111101011111110111110101110100010100000111111101111101011111010111010001110100010100000101000001000000011111110111110101111101011101000111010001010000010100000100000001111101011101000101000001000000010100000100000000000000000000000") port map( O =>C_31_S_4_out, I0 =>  C_31_S_4_L_0_out, I1 =>  C_31_S_4_L_1_out, I2 =>  C_31_S_4_L_2_out, I3 =>  C_31_S_4_L_3_out, I4 =>  C_31_S_4_L_4_out, I5 =>  C_31_S_4_L_5_out, I6 =>  C_31_S_4_L_6_out, I7 =>  C_31_S_4_L_7_out); 

C_31_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_31_out, I0 =>  C_31_S_0_out, I1 =>  C_31_S_1_out, I2 =>  C_31_S_2_out, I3 =>  C_31_S_3_out, I4 =>  C_31_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_32_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_32_S_0_out, I0 =>  C_32_S_0_L_0_out, I1 =>  C_32_S_0_L_1_out, I2 =>  C_32_S_0_L_2_out, I3 =>  C_32_S_0_L_3_out, I4 =>  C_32_S_0_L_4_out, I5 =>  C_32_S_0_L_5_out, I6 =>  C_32_S_0_L_6_out, I7 =>  C_32_S_0_L_7_out); 
C_32_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_32_S_1_out, I0 =>  C_32_S_1_L_0_out, I1 =>  C_32_S_1_L_1_out, I2 =>  C_32_S_1_L_2_out, I3 =>  C_32_S_1_L_3_out, I4 =>  C_32_S_1_L_4_out, I5 =>  C_32_S_1_L_5_out, I6 =>  C_32_S_1_L_6_out, I7 =>  C_32_S_1_L_7_out); 
C_32_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_32_S_2_out, I0 =>  C_32_S_2_L_0_out, I1 =>  C_32_S_2_L_1_out, I2 =>  C_32_S_2_L_2_out, I3 =>  C_32_S_2_L_3_out, I4 =>  C_32_S_2_L_4_out, I5 =>  C_32_S_2_L_5_out, I6 =>  C_32_S_2_L_6_out, I7 =>  C_32_S_2_L_7_out); 
C_32_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_32_S_3_out, I0 =>  C_32_S_3_L_0_out, I1 =>  C_32_S_3_L_1_out, I2 =>  C_32_S_3_L_2_out, I3 =>  C_32_S_3_L_3_out, I4 =>  C_32_S_3_L_4_out, I5 =>  C_32_S_3_L_5_out, I6 =>  C_32_S_3_L_6_out, I7 =>  C_32_S_3_L_7_out); 
C_32_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_32_S_4_out, I0 =>  C_32_S_4_L_0_out, I1 =>  C_32_S_4_L_1_out, I2 =>  C_32_S_4_L_2_out, I3 =>  C_32_S_4_L_3_out, I4 =>  C_32_S_4_L_4_out, I5 =>  C_32_S_4_L_5_out, I6 =>  C_32_S_4_L_6_out, I7 =>  C_32_S_4_L_7_out); 

C_32_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_32_out, I0 =>  C_32_S_0_out, I1 =>  C_32_S_1_out, I2 =>  C_32_S_2_out, I3 =>  C_32_S_3_out, I4 =>  C_32_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_33_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_33_S_0_out, I0 =>  C_33_S_0_L_0_out, I1 =>  C_33_S_0_L_1_out, I2 =>  C_33_S_0_L_2_out, I3 =>  C_33_S_0_L_3_out, I4 =>  C_33_S_0_L_4_out, I5 =>  C_33_S_0_L_5_out, I6 =>  C_33_S_0_L_6_out, I7 =>  C_33_S_0_L_7_out); 
C_33_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111110011111100100000001111100010000000100000000000000011111111111111101111111011100000111111101100000011000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_33_S_1_out, I0 =>  C_33_S_1_L_0_out, I1 =>  C_33_S_1_L_1_out, I2 =>  C_33_S_1_L_2_out, I3 =>  C_33_S_1_L_3_out, I4 =>  C_33_S_1_L_4_out, I5 =>  C_33_S_1_L_5_out, I6 =>  C_33_S_1_L_6_out, I7 =>  C_33_S_1_L_7_out); 
C_33_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_33_S_2_out, I0 =>  C_33_S_2_L_0_out, I1 =>  C_33_S_2_L_1_out, I2 =>  C_33_S_2_L_2_out, I3 =>  C_33_S_2_L_3_out, I4 =>  C_33_S_2_L_4_out, I5 =>  C_33_S_2_L_5_out, I6 =>  C_33_S_2_L_6_out, I7 =>  C_33_S_2_L_7_out); 
C_33_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_33_S_3_out, I0 =>  C_33_S_3_L_0_out, I1 =>  C_33_S_3_L_1_out, I2 =>  C_33_S_3_L_2_out, I3 =>  C_33_S_3_L_3_out, I4 =>  C_33_S_3_L_4_out, I5 =>  C_33_S_3_L_5_out, I6 =>  C_33_S_3_L_6_out, I7 =>  C_33_S_3_L_7_out); 
C_33_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111101011111110101000001111100010000000100000000000000011111111111111101111111011100000111110101000000010100000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_33_S_4_out, I0 =>  C_33_S_4_L_0_out, I1 =>  C_33_S_4_L_1_out, I2 =>  C_33_S_4_L_2_out, I3 =>  C_33_S_4_L_3_out, I4 =>  C_33_S_4_L_4_out, I5 =>  C_33_S_4_L_5_out, I6 =>  C_33_S_4_L_6_out, I7 =>  C_33_S_4_L_7_out); 

C_33_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_33_out, I0 =>  C_33_S_0_out, I1 =>  C_33_S_1_out, I2 =>  C_33_S_2_out, I3 =>  C_33_S_3_out, I4 =>  C_33_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_34_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_34_S_0_out, I0 =>  C_34_S_0_L_0_out, I1 =>  C_34_S_0_L_1_out, I2 =>  C_34_S_0_L_2_out, I3 =>  C_34_S_0_L_3_out, I4 =>  C_34_S_0_L_4_out, I5 =>  C_34_S_0_L_5_out, I6 =>  C_34_S_0_L_6_out, I7 =>  C_34_S_0_L_7_out); 
C_34_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111010100000001111111011101000100000000000000011111111111111101110100010000000111111101010000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_34_S_1_out, I0 =>  C_34_S_1_L_0_out, I1 =>  C_34_S_1_L_1_out, I2 =>  C_34_S_1_L_2_out, I3 =>  C_34_S_1_L_3_out, I4 =>  C_34_S_1_L_4_out, I5 =>  C_34_S_1_L_5_out, I6 =>  C_34_S_1_L_6_out, I7 =>  C_34_S_1_L_7_out); 
C_34_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111111110100011111110111010001110111010000000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001111111010001000111010001000000011101000000000001000000000000000") port map( O =>C_34_S_2_out, I0 =>  C_34_S_2_L_0_out, I1 =>  C_34_S_2_L_1_out, I2 =>  C_34_S_2_L_2_out, I3 =>  C_34_S_2_L_3_out, I4 =>  C_34_S_2_L_4_out, I5 =>  C_34_S_2_L_5_out, I6 =>  C_34_S_2_L_6_out, I7 =>  C_34_S_2_L_7_out); 
C_34_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101111111011111110111111101110100011101000111111101110100011101000100000001110100010000000100000001000000011111110111111101111111011101000111111101110100011101000100000001110100011101000100000001000000010000000100000001000000000000000") port map( O =>C_34_S_3_out, I0 =>  C_34_S_3_L_0_out, I1 =>  C_34_S_3_L_1_out, I2 =>  C_34_S_3_L_2_out, I3 =>  C_34_S_3_L_3_out, I4 =>  C_34_S_3_L_4_out, I5 =>  C_34_S_3_L_5_out, I6 =>  C_34_S_3_L_6_out, I7 =>  C_34_S_3_L_7_out); 
C_34_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101111111011101000111010001110100011101000100000001000000011111110111111101110100011101000111010001110100010000000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_34_S_4_out, I0 =>  C_34_S_4_L_0_out, I1 =>  C_34_S_4_L_1_out, I2 =>  C_34_S_4_L_2_out, I3 =>  C_34_S_4_L_3_out, I4 =>  C_34_S_4_L_4_out, I5 =>  C_34_S_4_L_5_out, I6 =>  C_34_S_4_L_6_out, I7 =>  C_34_S_4_L_7_out); 

C_34_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_34_out, I0 =>  C_34_S_0_out, I1 =>  C_34_S_1_out, I2 =>  C_34_S_2_out, I3 =>  C_34_S_3_out, I4 =>  C_34_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_35_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111011101110111011101000111111101110111011101010101010001110111010101000101010001000000011111110111010101110101010001000111010101010100010001000100000001110100010001000100010001000000010001000100000001000000000000000") port map( O =>C_35_S_0_out, I0 =>  C_35_S_0_L_0_out, I1 =>  C_35_S_0_L_1_out, I2 =>  C_35_S_0_L_2_out, I3 =>  C_35_S_0_L_3_out, I4 =>  C_35_S_0_L_4_out, I5 =>  C_35_S_0_L_5_out, I6 =>  C_35_S_0_L_6_out, I7 =>  C_35_S_0_L_7_out); 
C_35_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100011100000111111101110100011101000101000001110100011101000111000001000000011111110111110001110100011101000111110101110100011101000100000001111100011101000111010001000000011101000100000001000000000000000") port map( O =>C_35_S_1_out, I0 =>  C_35_S_1_L_0_out, I1 =>  C_35_S_1_L_1_out, I2 =>  C_35_S_1_L_2_out, I3 =>  C_35_S_1_L_3_out, I4 =>  C_35_S_1_L_4_out, I5 =>  C_35_S_1_L_5_out, I6 =>  C_35_S_1_L_6_out, I7 =>  C_35_S_1_L_7_out); 
C_35_S_2_inst : LUT8 generic map(INIT => "1111111011111000111111101110100011111110111010001111111011101000111111101110100011111110111010001111100011101000111010001000000011111110111010001110100011100000111010001000000011101000100000001110100010000000111010001000000011101000100000001110000010000000") port map( O =>C_35_S_2_out, I0 =>  C_35_S_2_L_0_out, I1 =>  C_35_S_2_L_1_out, I2 =>  C_35_S_2_L_2_out, I3 =>  C_35_S_2_L_3_out, I4 =>  C_35_S_2_L_4_out, I5 =>  C_35_S_2_L_5_out, I6 =>  C_35_S_2_L_6_out, I7 =>  C_35_S_2_L_7_out); 
C_35_S_3_inst : LUT8 generic map(INIT => "1111111011101000111111101110100011111110111010001111111011101000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001110100010000000111010001000000011101000100000001110100010000000") port map( O =>C_35_S_3_out, I0 =>  C_35_S_3_L_0_out, I1 =>  C_35_S_3_L_1_out, I2 =>  C_35_S_3_L_2_out, I3 =>  C_35_S_3_L_3_out, I4 =>  C_35_S_3_L_4_out, I5 =>  C_35_S_3_L_5_out, I6 =>  C_35_S_3_L_6_out, I7 =>  C_35_S_3_L_7_out); 
C_35_S_4_inst : LUT8 generic map(INIT => "1111111011101000111111101110100011111110111010001111111011101000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001110100010000000111010001000000011101000100000001110100010000000") port map( O =>C_35_S_4_out, I0 =>  C_35_S_4_L_0_out, I1 =>  C_35_S_4_L_1_out, I2 =>  C_35_S_4_L_2_out, I3 =>  C_35_S_4_L_3_out, I4 =>  C_35_S_4_L_4_out, I5 =>  C_35_S_4_L_5_out, I6 =>  C_35_S_4_L_6_out, I7 =>  C_35_S_4_L_7_out); 

C_35_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_35_out, I0 =>  C_35_S_0_out, I1 =>  C_35_S_1_out, I2 =>  C_35_S_2_out, I3 =>  C_35_S_3_out, I4 =>  C_35_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_36_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111111111011111110111010001110100010000000100000000000000011111111111111101111111011101000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_36_S_0_out, I0 =>  C_36_S_0_L_0_out, I1 =>  C_36_S_0_L_1_out, I2 =>  C_36_S_0_L_2_out, I3 =>  C_36_S_0_L_3_out, I4 =>  C_36_S_0_L_4_out, I5 =>  C_36_S_0_L_5_out, I6 =>  C_36_S_0_L_6_out, I7 =>  C_36_S_0_L_7_out); 
C_36_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_36_S_1_out, I0 =>  C_36_S_1_L_0_out, I1 =>  C_36_S_1_L_1_out, I2 =>  C_36_S_1_L_2_out, I3 =>  C_36_S_1_L_3_out, I4 =>  C_36_S_1_L_4_out, I5 =>  C_36_S_1_L_5_out, I6 =>  C_36_S_1_L_6_out, I7 =>  C_36_S_1_L_7_out); 
C_36_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111011101110111011001000111111111111111011101110110010001110111011001000100010001000000011111110111011101110110010001000111011001000100010000000000000001110110010001000100010000000000010000000000000000000000000000000") port map( O =>C_36_S_2_out, I0 =>  C_36_S_2_L_0_out, I1 =>  C_36_S_2_L_1_out, I2 =>  C_36_S_2_L_2_out, I3 =>  C_36_S_2_L_3_out, I4 =>  C_36_S_2_L_4_out, I5 =>  C_36_S_2_L_5_out, I6 =>  C_36_S_2_L_6_out, I7 =>  C_36_S_2_L_7_out); 
C_36_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111110111111101110100011101000111111101111111011101100111010001110100011101000100000001000000011111110111111101110100011101000111010001100100010000000100000001110100011101000100000001000000010000000000000000000000000000000") port map( O =>C_36_S_3_out, I0 =>  C_36_S_3_L_0_out, I1 =>  C_36_S_3_L_1_out, I2 =>  C_36_S_3_L_2_out, I3 =>  C_36_S_3_L_3_out, I4 =>  C_36_S_3_L_4_out, I5 =>  C_36_S_3_L_5_out, I6 =>  C_36_S_3_L_6_out, I7 =>  C_36_S_3_L_7_out); 
C_36_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111011101110100011101000111111101111111011101000111010001111111011101000111010001000000011111110111010001110100010000000111010001110100010000000100000001110100011101000100010001000000011101000100000001000000000000000") port map( O =>C_36_S_4_out, I0 =>  C_36_S_4_L_0_out, I1 =>  C_36_S_4_L_1_out, I2 =>  C_36_S_4_L_2_out, I3 =>  C_36_S_4_L_3_out, I4 =>  C_36_S_4_L_4_out, I5 =>  C_36_S_4_L_5_out, I6 =>  C_36_S_4_L_6_out, I7 =>  C_36_S_4_L_7_out); 

C_36_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_36_out, I0 =>  C_36_S_0_out, I1 =>  C_36_S_1_out, I2 =>  C_36_S_2_out, I3 =>  C_36_S_3_out, I4 =>  C_36_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_37_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010001110100010000000111111101110101011101010111010001110100010101000100010001000000011111110111011101110101011101000111010001010100010101000100000001111111011101000111010001000000010101000100000001000000000000000") port map( O =>C_37_S_0_out, I0 =>  C_37_S_0_L_0_out, I1 =>  C_37_S_0_L_1_out, I2 =>  C_37_S_0_L_2_out, I3 =>  C_37_S_0_L_3_out, I4 =>  C_37_S_0_L_4_out, I5 =>  C_37_S_0_L_5_out, I6 =>  C_37_S_0_L_6_out, I7 =>  C_37_S_0_L_7_out); 
C_37_S_1_inst : LUT8 generic map(INIT => "1111111011111110111111101111111011111110111010001110100011101000111111101110100011101010111010001110100011101000111010001000000011111110111010001110100011101000111010001010100011101000100000001110100011101000111010001000000010000000100000001000000010000000") port map( O =>C_37_S_1_out, I0 =>  C_37_S_1_L_0_out, I1 =>  C_37_S_1_L_1_out, I2 =>  C_37_S_1_L_2_out, I3 =>  C_37_S_1_L_3_out, I4 =>  C_37_S_1_L_4_out, I5 =>  C_37_S_1_L_5_out, I6 =>  C_37_S_1_L_6_out, I7 =>  C_37_S_1_L_7_out); 
C_37_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111011101110100011101000111111101110111011101000111010001110111011101000111010001000000011111110111010001110100010001000111010001110100010001000100000001110100011101000100010001000000011101000100000001000000000000000") port map( O =>C_37_S_2_out, I0 =>  C_37_S_2_L_0_out, I1 =>  C_37_S_2_L_1_out, I2 =>  C_37_S_2_L_2_out, I3 =>  C_37_S_2_L_3_out, I4 =>  C_37_S_2_L_4_out, I5 =>  C_37_S_2_L_5_out, I6 =>  C_37_S_2_L_6_out, I7 =>  C_37_S_2_L_7_out); 
C_37_S_3_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111010111010001110100011101000111111101111101011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100010100000100000001110100011101000111010001010000011101000100000001000000010000000") port map( O =>C_37_S_3_out, I0 =>  C_37_S_3_L_0_out, I1 =>  C_37_S_3_L_1_out, I2 =>  C_37_S_3_L_2_out, I3 =>  C_37_S_3_L_3_out, I4 =>  C_37_S_3_L_4_out, I5 =>  C_37_S_3_L_5_out, I6 =>  C_37_S_3_L_6_out, I7 =>  C_37_S_3_L_7_out); 
C_37_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010101110100011101000111111101110100011101000101010001110100011101000101010001000000011111110111010101110100011101000111010101110100011101000100000001110100011101000101010001000000011101000100000001000000000000000") port map( O =>C_37_S_4_out, I0 =>  C_37_S_4_L_0_out, I1 =>  C_37_S_4_L_1_out, I2 =>  C_37_S_4_L_2_out, I3 =>  C_37_S_4_L_3_out, I4 =>  C_37_S_4_L_4_out, I5 =>  C_37_S_4_L_5_out, I6 =>  C_37_S_4_L_6_out, I7 =>  C_37_S_4_L_7_out); 

C_37_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_37_out, I0 =>  C_37_S_0_out, I1 =>  C_37_S_1_out, I2 =>  C_37_S_2_out, I3 =>  C_37_S_3_out, I4 =>  C_37_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_38_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111101011111111111110101111101010100000111111111111101011111010101000001111101010100000101000000000000011111111111110101111101010100000111110101010000010100000000000001111101010100000101000000000000010100000000000000000000000000000") port map( O =>C_38_S_0_out, I0 =>  C_38_S_0_L_0_out, I1 =>  C_38_S_0_L_1_out, I2 =>  C_38_S_0_L_2_out, I3 =>  C_38_S_0_L_3_out, I4 =>  C_38_S_0_L_4_out, I5 =>  C_38_S_0_L_5_out, I6 =>  C_38_S_0_L_6_out, I7 =>  C_38_S_0_L_7_out); 
C_38_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111110111010001111111011100000111010000000000011111111111010001111100010000000111010001000000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_38_S_1_out, I0 =>  C_38_S_1_L_0_out, I1 =>  C_38_S_1_L_1_out, I2 =>  C_38_S_1_L_2_out, I3 =>  C_38_S_1_L_3_out, I4 =>  C_38_S_1_L_4_out, I5 =>  C_38_S_1_L_5_out, I6 =>  C_38_S_1_L_6_out, I7 =>  C_38_S_1_L_7_out); 
C_38_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111101111100011111110111110001110100010000000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001111111011101000111000001000000011100000100000000000000000000000") port map( O =>C_38_S_2_out, I0 =>  C_38_S_2_L_0_out, I1 =>  C_38_S_2_L_1_out, I2 =>  C_38_S_2_L_2_out, I3 =>  C_38_S_2_L_3_out, I4 =>  C_38_S_2_L_4_out, I5 =>  C_38_S_2_L_5_out, I6 =>  C_38_S_2_L_6_out, I7 =>  C_38_S_2_L_7_out); 
C_38_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111110111010001111111011101000111010001000000011111110111010001110100010000000111010001000000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_38_S_3_out, I0 =>  C_38_S_3_L_0_out, I1 =>  C_38_S_3_L_1_out, I2 =>  C_38_S_3_L_2_out, I3 =>  C_38_S_3_L_3_out, I4 =>  C_38_S_3_L_4_out, I5 =>  C_38_S_3_L_5_out, I6 =>  C_38_S_3_L_6_out, I7 =>  C_38_S_3_L_7_out); 
C_38_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010000000000011111111111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_38_S_4_out, I0 =>  C_38_S_4_L_0_out, I1 =>  C_38_S_4_L_1_out, I2 =>  C_38_S_4_L_2_out, I3 =>  C_38_S_4_L_3_out, I4 =>  C_38_S_4_L_4_out, I5 =>  C_38_S_4_L_5_out, I6 =>  C_38_S_4_L_6_out, I7 =>  C_38_S_4_L_7_out); 

C_38_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_38_out, I0 =>  C_38_S_0_out, I1 =>  C_38_S_1_out, I2 =>  C_38_S_2_out, I3 =>  C_38_S_3_out, I4 =>  C_38_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_39_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100011100000111111101110100011101000111000001110100011101000111000001000000011111110111110001110100011101000111110001110100011101000100000001111100011101000111010001000000011101000100000001000000000000000") port map( O =>C_39_S_0_out, I0 =>  C_39_S_0_L_0_out, I1 =>  C_39_S_0_L_1_out, I2 =>  C_39_S_0_L_2_out, I3 =>  C_39_S_0_L_3_out, I4 =>  C_39_S_0_L_4_out, I5 =>  C_39_S_0_L_5_out, I6 =>  C_39_S_0_L_6_out, I7 =>  C_39_S_0_L_7_out); 
C_39_S_1_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_39_S_1_out, I0 =>  C_39_S_1_L_0_out, I1 =>  C_39_S_1_L_1_out, I2 =>  C_39_S_1_L_2_out, I3 =>  C_39_S_1_L_3_out, I4 =>  C_39_S_1_L_4_out, I5 =>  C_39_S_1_L_5_out, I6 =>  C_39_S_1_L_6_out, I7 =>  C_39_S_1_L_7_out); 
C_39_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110111010101000111111101110100011101000100010001110101010101000101010001000000011111110111010101110101010101000111011101110100011101000100000001110101010001000101010001000000010101000100000001000000000000000") port map( O =>C_39_S_2_out, I0 =>  C_39_S_2_L_0_out, I1 =>  C_39_S_2_L_1_out, I2 =>  C_39_S_2_L_2_out, I3 =>  C_39_S_2_L_3_out, I4 =>  C_39_S_2_L_4_out, I5 =>  C_39_S_2_L_5_out, I6 =>  C_39_S_2_L_6_out, I7 =>  C_39_S_2_L_7_out); 
C_39_S_3_inst : LUT8 generic map(INIT => "1111111011111000111111101110100011111110111010001111101011101000111111101110100011111000101000001111101011101000111010001000000011111110111010001110100010100000111110101110000011101000100000001110100010100000111010001000000011101000100000001110000010000000") port map( O =>C_39_S_3_out, I0 =>  C_39_S_3_L_0_out, I1 =>  C_39_S_3_L_1_out, I2 =>  C_39_S_3_L_2_out, I3 =>  C_39_S_3_L_3_out, I4 =>  C_39_S_3_L_4_out, I5 =>  C_39_S_3_L_5_out, I6 =>  C_39_S_3_L_6_out, I7 =>  C_39_S_3_L_7_out); 
C_39_S_4_inst : LUT8 generic map(INIT => "1111111011111110111110101110100011111110111010001110100011101000111111101110100011101000111010001111100011101000111010001000000011111110111010001110100011100000111010001110100011101000100000001110100011101000111010001000000011101000101000001000000010000000") port map( O =>C_39_S_4_out, I0 =>  C_39_S_4_L_0_out, I1 =>  C_39_S_4_L_1_out, I2 =>  C_39_S_4_L_2_out, I3 =>  C_39_S_4_L_3_out, I4 =>  C_39_S_4_L_4_out, I5 =>  C_39_S_4_L_5_out, I6 =>  C_39_S_4_L_6_out, I7 =>  C_39_S_4_L_7_out); 

C_39_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_39_out, I0 =>  C_39_S_0_out, I1 =>  C_39_S_1_out, I2 =>  C_39_S_2_out, I3 =>  C_39_S_3_out, I4 =>  C_39_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_40_S_0_inst : LUT8 generic map(INIT => "1111111011101110111011101110111011101110111010101110101011101000111011101110101011101000111010001110100010101000101010001000100011101110111010101110101011101000111010001110100010101000100010001110100010101000101010001000100010001000100010001000100010000000") port map( O =>C_40_S_0_out, I0 =>  C_40_S_0_L_0_out, I1 =>  C_40_S_0_L_1_out, I2 =>  C_40_S_0_L_2_out, I3 =>  C_40_S_0_L_3_out, I4 =>  C_40_S_0_L_4_out, I5 =>  C_40_S_0_L_5_out, I6 =>  C_40_S_0_L_6_out, I7 =>  C_40_S_0_L_7_out); 
C_40_S_1_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010001110100010101000111011101110101011101010111010001110100010101000101010001000100011101110111010101110101011101000111010001010100010101000100010001110101011101000111010001000100010101000100010001000100010000000") port map( O =>C_40_S_1_out, I0 =>  C_40_S_1_L_0_out, I1 =>  C_40_S_1_L_1_out, I2 =>  C_40_S_1_L_2_out, I3 =>  C_40_S_1_L_3_out, I4 =>  C_40_S_1_L_4_out, I5 =>  C_40_S_1_L_5_out, I6 =>  C_40_S_1_L_6_out, I7 =>  C_40_S_1_L_7_out); 
C_40_S_2_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010101110101010101000111011101110101011101010101010001110101010101000111010001000100011101110111010001110101010101000111010101010100010101000100010001110101010101000101010001000100011101000100010001000100010000000") port map( O =>C_40_S_2_out, I0 =>  C_40_S_2_L_0_out, I1 =>  C_40_S_2_L_1_out, I2 =>  C_40_S_2_L_2_out, I3 =>  C_40_S_2_L_3_out, I4 =>  C_40_S_2_L_4_out, I5 =>  C_40_S_2_L_5_out, I6 =>  C_40_S_2_L_6_out, I7 =>  C_40_S_2_L_7_out); 
C_40_S_3_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_40_S_3_out, I0 =>  C_40_S_3_L_0_out, I1 =>  C_40_S_3_L_1_out, I2 =>  C_40_S_3_L_2_out, I3 =>  C_40_S_3_L_3_out, I4 =>  C_40_S_3_L_4_out, I5 =>  C_40_S_3_L_5_out, I6 =>  C_40_S_3_L_6_out, I7 =>  C_40_S_3_L_7_out); 
C_40_S_4_inst : LUT8 generic map(INIT => "1111111011101010111110101110100011111010111010001110101010101000111111101110101011101010101010001110101010101000101010001010000011111010111010101110101010101000111010101010100010101000100000001110101010101000111010001010000011101000101000001010100010000000") port map( O =>C_40_S_4_out, I0 =>  C_40_S_4_L_0_out, I1 =>  C_40_S_4_L_1_out, I2 =>  C_40_S_4_L_2_out, I3 =>  C_40_S_4_L_3_out, I4 =>  C_40_S_4_L_4_out, I5 =>  C_40_S_4_L_5_out, I6 =>  C_40_S_4_L_6_out, I7 =>  C_40_S_4_L_7_out); 

C_40_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_40_out, I0 =>  C_40_S_0_out, I1 =>  C_40_S_1_out, I2 =>  C_40_S_2_out, I3 =>  C_40_S_3_out, I4 =>  C_40_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_41_S_0_inst : LUT8 generic map(INIT => "1110111011101110111011101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100010001000100010001000") port map( O =>C_41_S_0_out, I0 =>  C_41_S_0_L_0_out, I1 =>  C_41_S_0_L_1_out, I2 =>  C_41_S_0_L_2_out, I3 =>  C_41_S_0_L_3_out, I4 =>  C_41_S_0_L_4_out, I5 =>  C_41_S_0_L_5_out, I6 =>  C_41_S_0_L_6_out, I7 =>  C_41_S_0_L_7_out); 
C_41_S_1_inst : LUT8 generic map(INIT => "1111111111111110111011101110100011101110111010001110100010001000111111101110111011101000111010001110100011101000100010001000000011111110111011101110100011101000111010001110100010001000100000001110111011101000111010001000100011101000100010001000000000000000") port map( O =>C_41_S_1_out, I0 =>  C_41_S_1_L_0_out, I1 =>  C_41_S_1_L_1_out, I2 =>  C_41_S_1_L_2_out, I3 =>  C_41_S_1_L_3_out, I4 =>  C_41_S_1_L_4_out, I5 =>  C_41_S_1_L_5_out, I6 =>  C_41_S_1_L_6_out, I7 =>  C_41_S_1_L_7_out); 
C_41_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010001110100010101000111111101110101011101010111010001110100010101000101010001000000011111110111010101110101011101000111010001010100010101000100000001110101011101000111010001000000010101000100000001000000000000000") port map( O =>C_41_S_2_out, I0 =>  C_41_S_2_L_0_out, I1 =>  C_41_S_2_L_1_out, I2 =>  C_41_S_2_L_2_out, I3 =>  C_41_S_2_L_3_out, I4 =>  C_41_S_2_L_4_out, I5 =>  C_41_S_2_L_5_out, I6 =>  C_41_S_2_L_6_out, I7 =>  C_41_S_2_L_7_out); 
C_41_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101010101011111111111010101110101010100000111111101010101010101010100000001110101010101000101010000000000011111111111010101110101010101000111111101010101010101010100000001111101010101000101010000000000010101010100000001000000000000000") port map( O =>C_41_S_3_out, I0 =>  C_41_S_3_L_0_out, I1 =>  C_41_S_3_L_1_out, I2 =>  C_41_S_3_L_2_out, I3 =>  C_41_S_3_L_3_out, I4 =>  C_41_S_3_L_4_out, I5 =>  C_41_S_3_L_5_out, I6 =>  C_41_S_3_L_6_out, I7 =>  C_41_S_3_L_7_out); 
C_41_S_4_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_41_S_4_out, I0 =>  C_41_S_4_L_0_out, I1 =>  C_41_S_4_L_1_out, I2 =>  C_41_S_4_L_2_out, I3 =>  C_41_S_4_L_3_out, I4 =>  C_41_S_4_L_4_out, I5 =>  C_41_S_4_L_5_out, I6 =>  C_41_S_4_L_6_out, I7 =>  C_41_S_4_L_7_out); 

C_41_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_41_out, I0 =>  C_41_S_0_out, I1 =>  C_41_S_1_out, I2 =>  C_41_S_2_out, I3 =>  C_41_S_3_out, I4 =>  C_41_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_42_S_0_inst : LUT8 generic map(INIT => "1111111011111110111011101110101011101110111011101110100010101000111011101110111011101000101010001110101011101000101010001000100011101110111010101110100010101000111010101110100010001000100010001110101011101000100010001000100010101000100010001000000010000000") port map( O =>C_42_S_0_out, I0 =>  C_42_S_0_L_0_out, I1 =>  C_42_S_0_L_1_out, I2 =>  C_42_S_0_L_2_out, I3 =>  C_42_S_0_L_3_out, I4 =>  C_42_S_0_L_4_out, I5 =>  C_42_S_0_L_5_out, I6 =>  C_42_S_0_L_6_out, I7 =>  C_42_S_0_L_7_out); 
C_42_S_1_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010001110111010001000111011101110100011101110100010001110100010001000100010001000100011101110111011101110111011101000111011101000100011101000100010001110111010001000111010001000100010101000100010001000100010000000") port map( O =>C_42_S_1_out, I0 =>  C_42_S_1_L_0_out, I1 =>  C_42_S_1_L_1_out, I2 =>  C_42_S_1_L_2_out, I3 =>  C_42_S_1_L_3_out, I4 =>  C_42_S_1_L_4_out, I5 =>  C_42_S_1_L_5_out, I6 =>  C_42_S_1_L_6_out, I7 =>  C_42_S_1_L_7_out); 
C_42_S_2_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010001110101010101000111011101110100011101010101010001110101011101000111010001000100011101110111010001110100010101000111010101010100011101000100010001110101010101000111010001000100011101000100010001000100010000000") port map( O =>C_42_S_2_out, I0 =>  C_42_S_2_L_0_out, I1 =>  C_42_S_2_L_1_out, I2 =>  C_42_S_2_L_2_out, I3 =>  C_42_S_2_L_3_out, I4 =>  C_42_S_2_L_4_out, I5 =>  C_42_S_2_L_5_out, I6 =>  C_42_S_2_L_6_out, I7 =>  C_42_S_2_L_7_out); 
C_42_S_3_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010101110100010101000111011101110101011101000101010001110101010101000101010001000100011101110111010101110101010101000111010101110100010101000100010001110101011101000101010001000100011101000100010001000100010000000") port map( O =>C_42_S_3_out, I0 =>  C_42_S_3_L_0_out, I1 =>  C_42_S_3_L_1_out, I2 =>  C_42_S_3_L_2_out, I3 =>  C_42_S_3_L_3_out, I4 =>  C_42_S_3_L_4_out, I5 =>  C_42_S_3_L_5_out, I6 =>  C_42_S_3_L_6_out, I7 =>  C_42_S_3_L_7_out); 
C_42_S_4_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010101110100010101000111011101110101011101000101010001110101011101000101010001000100011101110111010101110100010101000111010101110100010101000100010001110101011101000101010001000100011101000100010001000100010000000") port map( O =>C_42_S_4_out, I0 =>  C_42_S_4_L_0_out, I1 =>  C_42_S_4_L_1_out, I2 =>  C_42_S_4_L_2_out, I3 =>  C_42_S_4_L_3_out, I4 =>  C_42_S_4_L_4_out, I5 =>  C_42_S_4_L_5_out, I6 =>  C_42_S_4_L_6_out, I7 =>  C_42_S_4_L_7_out); 

C_42_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_42_out, I0 =>  C_42_S_0_out, I1 =>  C_42_S_1_out, I2 =>  C_42_S_2_out, I3 =>  C_42_S_3_out, I4 =>  C_42_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_43_S_0_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100011101000100010001000100010000000") port map( O =>C_43_S_0_out, I0 =>  C_43_S_0_L_0_out, I1 =>  C_43_S_0_L_1_out, I2 =>  C_43_S_0_L_2_out, I3 =>  C_43_S_0_L_3_out, I4 =>  C_43_S_0_L_4_out, I5 =>  C_43_S_0_L_5_out, I6 =>  C_43_S_0_L_6_out, I7 =>  C_43_S_0_L_7_out); 
C_43_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101110111010101110101010101000111010101010101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101010101010001110101010101000101010001000100010101010101010001010100010000000") port map( O =>C_43_S_1_out, I0 =>  C_43_S_1_L_0_out, I1 =>  C_43_S_1_L_1_out, I2 =>  C_43_S_1_L_2_out, I3 =>  C_43_S_1_L_3_out, I4 =>  C_43_S_1_L_4_out, I5 =>  C_43_S_1_L_5_out, I6 =>  C_43_S_1_L_6_out, I7 =>  C_43_S_1_L_7_out); 
C_43_S_2_inst : LUT8 generic map(INIT => "1111111011111110111111101110101011101010111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001010100010101000100000001000000010000000") port map( O =>C_43_S_2_out, I0 =>  C_43_S_2_L_0_out, I1 =>  C_43_S_2_L_1_out, I2 =>  C_43_S_2_L_2_out, I3 =>  C_43_S_2_L_3_out, I4 =>  C_43_S_2_L_4_out, I5 =>  C_43_S_2_L_5_out, I6 =>  C_43_S_2_L_6_out, I7 =>  C_43_S_2_L_7_out); 
C_43_S_3_inst : LUT8 generic map(INIT => "1111111011101110111111101110101011101010101010101110101010101010111010101010101011101010101010101010101010101000101010101010100011101010101010101110101010101010101010101010100010101010101010001010101010101000101010101010100010101000100000001000100010000000") port map( O =>C_43_S_3_out, I0 =>  C_43_S_3_L_0_out, I1 =>  C_43_S_3_L_1_out, I2 =>  C_43_S_3_L_2_out, I3 =>  C_43_S_3_L_3_out, I4 =>  C_43_S_3_L_4_out, I5 =>  C_43_S_3_L_5_out, I6 =>  C_43_S_3_L_6_out, I7 =>  C_43_S_3_L_7_out); 
C_43_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001111110011000000111111111111110011111110111010001111110011101000111010001000000011111110111010001110100011000000111010001000000011000000000000001111110011000000111010001000000011101000100000001000000000000000") port map( O =>C_43_S_4_out, I0 =>  C_43_S_4_L_0_out, I1 =>  C_43_S_4_L_1_out, I2 =>  C_43_S_4_L_2_out, I3 =>  C_43_S_4_L_3_out, I4 =>  C_43_S_4_L_4_out, I5 =>  C_43_S_4_L_5_out, I6 =>  C_43_S_4_L_6_out, I7 =>  C_43_S_4_L_7_out); 

C_43_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_43_out, I0 =>  C_43_S_0_out, I1 =>  C_43_S_1_out, I2 =>  C_43_S_2_out, I3 =>  C_43_S_3_out, I4 =>  C_43_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_44_S_0_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011111110111010101110101011101000111011101110100011101000100010001110101011101000111010001000100011101110111010001110100010101000111011101110100011101000100010001110100010101000101010001000000011101000100010001000100010000000") port map( O =>C_44_S_0_out, I0 =>  C_44_S_0_L_0_out, I1 =>  C_44_S_0_L_1_out, I2 =>  C_44_S_0_L_2_out, I3 =>  C_44_S_0_L_3_out, I4 =>  C_44_S_0_L_4_out, I5 =>  C_44_S_0_L_5_out, I6 =>  C_44_S_0_L_6_out, I7 =>  C_44_S_0_L_7_out); 
C_44_S_1_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010001110101010001000111011101110100011101110100010001110100010001000101010001000100011101110111010101110111011101000111011101000100011101000100010001110111010101000111010001000100011101000100010001000100010000000") port map( O =>C_44_S_1_out, I0 =>  C_44_S_1_L_0_out, I1 =>  C_44_S_1_L_1_out, I2 =>  C_44_S_1_L_2_out, I3 =>  C_44_S_1_L_3_out, I4 =>  C_44_S_1_L_4_out, I5 =>  C_44_S_1_L_5_out, I6 =>  C_44_S_1_L_6_out, I7 =>  C_44_S_1_L_7_out); 
C_44_S_2_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_44_S_2_out, I0 =>  C_44_S_2_L_0_out, I1 =>  C_44_S_2_L_1_out, I2 =>  C_44_S_2_L_2_out, I3 =>  C_44_S_2_L_3_out, I4 =>  C_44_S_2_L_4_out, I5 =>  C_44_S_2_L_5_out, I6 =>  C_44_S_2_L_6_out, I7 =>  C_44_S_2_L_7_out); 
C_44_S_3_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010001110101010101000111011101110101011101010111010001110100010001000101010001000100011101110111010101110111011101000111010001010100010101000100010001110101010101000111010001000100010101000100010001000100010000000") port map( O =>C_44_S_3_out, I0 =>  C_44_S_3_L_0_out, I1 =>  C_44_S_3_L_1_out, I2 =>  C_44_S_3_L_2_out, I3 =>  C_44_S_3_L_3_out, I4 =>  C_44_S_3_L_4_out, I5 =>  C_44_S_3_L_5_out, I6 =>  C_44_S_3_L_6_out, I7 =>  C_44_S_3_L_7_out); 
C_44_S_4_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100010001000100010000000") port map( O =>C_44_S_4_out, I0 =>  C_44_S_4_L_0_out, I1 =>  C_44_S_4_L_1_out, I2 =>  C_44_S_4_L_2_out, I3 =>  C_44_S_4_L_3_out, I4 =>  C_44_S_4_L_4_out, I5 =>  C_44_S_4_L_5_out, I6 =>  C_44_S_4_L_6_out, I7 =>  C_44_S_4_L_7_out); 

C_44_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_44_out, I0 =>  C_44_S_0_out, I1 =>  C_44_S_1_out, I2 =>  C_44_S_2_out, I3 =>  C_44_S_3_out, I4 =>  C_44_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_45_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101110101010101010101010101000111011101010101010101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010101010101010100010001110101010101010101010101000100010101010101010001010100010001000") port map( O =>C_45_S_0_out, I0 =>  C_45_S_0_L_0_out, I1 =>  C_45_S_0_L_1_out, I2 =>  C_45_S_0_L_2_out, I3 =>  C_45_S_0_L_3_out, I4 =>  C_45_S_0_L_4_out, I5 =>  C_45_S_0_L_5_out, I6 =>  C_45_S_0_L_6_out, I7 =>  C_45_S_0_L_7_out); 
C_45_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101110101010101000111010101010101011101010101010001110101010101000101010101010000011111010101010101110101010101000111010101010100010101010101010001110101010101000101010101010100010101010101010001010100010000000") port map( O =>C_45_S_1_out, I0 =>  C_45_S_1_L_0_out, I1 =>  C_45_S_1_L_1_out, I2 =>  C_45_S_1_L_2_out, I3 =>  C_45_S_1_L_3_out, I4 =>  C_45_S_1_L_4_out, I5 =>  C_45_S_1_L_5_out, I6 =>  C_45_S_1_L_6_out, I7 =>  C_45_S_1_L_7_out); 
C_45_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011101110111010101110101010101000111111101110111011101110111010001110101010101000101010001000000011111110111010101110101010101000111010001000100010001000100000001110101010101000101010001000100010001000100000001000000000000000") port map( O =>C_45_S_2_out, I0 =>  C_45_S_2_L_0_out, I1 =>  C_45_S_2_L_1_out, I2 =>  C_45_S_2_L_2_out, I3 =>  C_45_S_2_L_3_out, I4 =>  C_45_S_2_L_4_out, I5 =>  C_45_S_2_L_5_out, I6 =>  C_45_S_2_L_6_out, I7 =>  C_45_S_2_L_7_out); 
C_45_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111110110011111111111011001110110010000000111111111110111011111110100010001110111010000000110010000000000011111111111011001111111010001000111011101000000010001000000000001111111011001000110010000000000011001000000000000000000000000000") port map( O =>C_45_S_3_out, I0 =>  C_45_S_3_L_0_out, I1 =>  C_45_S_3_L_1_out, I2 =>  C_45_S_3_L_2_out, I3 =>  C_45_S_3_L_3_out, I4 =>  C_45_S_3_L_4_out, I5 =>  C_45_S_3_L_5_out, I6 =>  C_45_S_3_L_6_out, I7 =>  C_45_S_3_L_7_out); 
C_45_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101111111011111110111110101110100011101000111111101110100011101000111010001110100010100000100000001000000011111110111111101111101011101000111010001110100011101000100000001110100011101000101000001000000010000000100000001000000000000000") port map( O =>C_45_S_4_out, I0 =>  C_45_S_4_L_0_out, I1 =>  C_45_S_4_L_1_out, I2 =>  C_45_S_4_L_2_out, I3 =>  C_45_S_4_L_3_out, I4 =>  C_45_S_4_L_4_out, I5 =>  C_45_S_4_L_5_out, I6 =>  C_45_S_4_L_6_out, I7 =>  C_45_S_4_L_7_out); 

C_45_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_45_out, I0 =>  C_45_S_0_out, I1 =>  C_45_S_1_out, I2 =>  C_45_S_2_out, I3 =>  C_45_S_3_out, I4 =>  C_45_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_46_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010101110100010101000111111101110101011101000101010001110101011101000101010001000000011111110111010101110100010101000111010101110100010101000100000001110101011101000101010001000000011101000100000001000000000000000") port map( O =>C_46_S_0_out, I0 =>  C_46_S_0_L_0_out, I1 =>  C_46_S_0_L_1_out, I2 =>  C_46_S_0_L_2_out, I3 =>  C_46_S_0_L_3_out, I4 =>  C_46_S_0_L_4_out, I5 =>  C_46_S_0_L_5_out, I6 =>  C_46_S_0_L_6_out, I7 =>  C_46_S_0_L_7_out); 
C_46_S_1_inst : LUT8 generic map(INIT => "1111111111111110111011101110101011111110111011101110100010101000111111101110101011101000100010001110100010101000100010001000000011111110111011101110101011101000111011101110100010101000100000001110101011101000100010001000000010101000100010001000000000000000") port map( O =>C_46_S_1_out, I0 =>  C_46_S_1_L_0_out, I1 =>  C_46_S_1_L_1_out, I2 =>  C_46_S_1_L_2_out, I3 =>  C_46_S_1_L_3_out, I4 =>  C_46_S_1_L_4_out, I5 =>  C_46_S_1_L_5_out, I6 =>  C_46_S_1_L_6_out, I7 =>  C_46_S_1_L_7_out); 
C_46_S_2_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111011101110111010001000111011101110111011101110100010001110111011101000111010001000100011101110111010001110100010001000111011101000100010001000100010001110111010001000100010001000100011101000100010001000100010000000") port map( O =>C_46_S_2_out, I0 =>  C_46_S_2_L_0_out, I1 =>  C_46_S_2_L_1_out, I2 =>  C_46_S_2_L_2_out, I3 =>  C_46_S_2_L_3_out, I4 =>  C_46_S_2_L_4_out, I5 =>  C_46_S_2_L_5_out, I6 =>  C_46_S_2_L_6_out, I7 =>  C_46_S_2_L_7_out); 
C_46_S_3_inst : LUT8 generic map(INIT => "1111111011111110111011101110111011101110111011101110111011101000111011101110101011101000101010001110100010101000100010001000100011101110111011101110101011101000111010101110100010101000100010001110100010001000100010001000100010001000100010001000000010000000") port map( O =>C_46_S_3_out, I0 =>  C_46_S_3_L_0_out, I1 =>  C_46_S_3_L_1_out, I2 =>  C_46_S_3_L_2_out, I3 =>  C_46_S_3_L_3_out, I4 =>  C_46_S_3_L_4_out, I5 =>  C_46_S_3_L_5_out, I6 =>  C_46_S_3_L_6_out, I7 =>  C_46_S_3_L_7_out); 
C_46_S_4_inst : LUT8 generic map(INIT => "1111111011101110111011101110111011101110111010101110100010001000111011101110101011101000100010001110100010001000100010001000000011111110111011101110111011101000111011101110100010101000100010001110111011101000101010001000100010001000100010001000100010000000") port map( O =>C_46_S_4_out, I0 =>  C_46_S_4_L_0_out, I1 =>  C_46_S_4_L_1_out, I2 =>  C_46_S_4_L_2_out, I3 =>  C_46_S_4_L_3_out, I4 =>  C_46_S_4_L_4_out, I5 =>  C_46_S_4_L_5_out, I6 =>  C_46_S_4_L_6_out, I7 =>  C_46_S_4_L_7_out); 

C_46_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_46_out, I0 =>  C_46_S_0_out, I1 =>  C_46_S_1_out, I2 =>  C_46_S_2_out, I3 =>  C_46_S_3_out, I4 =>  C_46_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_47_S_0_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101110111010101110100010101000111011101110101011101000101010001110100010101000101010001000100011101110111010101110101011101000111010101110100010101000100010001110101011101000101010001000100010101000100010001000100010000000") port map( O =>C_47_S_0_out, I0 =>  C_47_S_0_L_0_out, I1 =>  C_47_S_0_L_1_out, I2 =>  C_47_S_0_L_2_out, I3 =>  C_47_S_0_L_3_out, I4 =>  C_47_S_0_L_4_out, I5 =>  C_47_S_0_L_5_out, I6 =>  C_47_S_0_L_6_out, I7 =>  C_47_S_0_L_7_out); 
C_47_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101000111110101110101011101010101010101110101010101010101010101010000011111010101010101010101010101000101010101010100010101000101000001110101010101010101010101010100010101010101010001010100010000000") port map( O =>C_47_S_1_out, I0 =>  C_47_S_1_L_0_out, I1 =>  C_47_S_1_L_1_out, I2 =>  C_47_S_1_L_2_out, I3 =>  C_47_S_1_L_3_out, I4 =>  C_47_S_1_L_4_out, I5 =>  C_47_S_1_L_5_out, I6 =>  C_47_S_1_L_6_out, I7 =>  C_47_S_1_L_7_out); 
C_47_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111110111011101110111010001110100010001000100000000000000011111111111111101110111011101000111010001000100010001000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_47_S_2_out, I0 =>  C_47_S_2_L_0_out, I1 =>  C_47_S_2_L_1_out, I2 =>  C_47_S_2_L_2_out, I3 =>  C_47_S_2_L_3_out, I4 =>  C_47_S_2_L_4_out, I5 =>  C_47_S_2_L_5_out, I6 =>  C_47_S_2_L_6_out, I7 =>  C_47_S_2_L_7_out); 
C_47_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111101110111011111111111111101111111011101000111111111111111011101000100000001111111011101000110010001000000011111110111011001110100010000000111111101110100010000000000000001110100010000000100000000000000010001000100000000000000000000000") port map( O =>C_47_S_3_out, I0 =>  C_47_S_3_L_0_out, I1 =>  C_47_S_3_L_1_out, I2 =>  C_47_S_3_L_2_out, I3 =>  C_47_S_3_L_3_out, I4 =>  C_47_S_3_L_4_out, I5 =>  C_47_S_3_L_5_out, I6 =>  C_47_S_3_L_6_out, I7 =>  C_47_S_3_L_7_out); 
C_47_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010001110101010001000111111101110111011101110111010001110111011101000111010001000000011111110111010001110100010001000111010001000100010001000100000001110111010101000111010001000000010101000100000001000000000000000") port map( O =>C_47_S_4_out, I0 =>  C_47_S_4_L_0_out, I1 =>  C_47_S_4_L_1_out, I2 =>  C_47_S_4_L_2_out, I3 =>  C_47_S_4_L_3_out, I4 =>  C_47_S_4_L_4_out, I5 =>  C_47_S_4_L_5_out, I6 =>  C_47_S_4_L_6_out, I7 =>  C_47_S_4_L_7_out); 

C_47_inst : LUT8 generic map(INIT => "1111101011101000111010001010000011111010111010001110100010100000111110101110100011101000101000001111101011101000111010001010000011111010111010001110100010100000111110101110100011101000101000001111101011101000111010001010000011111010111010001110100010100000") port map( O =>C_47_out, I0 =>  C_47_S_0_out, I1 =>  C_47_S_1_out, I2 =>  C_47_S_2_out, I3 =>  C_47_S_3_out, I4 =>  C_47_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_48_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101010101010101010101010101000111010101010101011101010101010101010101010101000101010001010100011101010111010101110101010101010101010101010100010101010101010001110101010101010101010101010100010101010101010001010100010001000") port map( O =>C_48_S_0_out, I0 =>  C_48_S_0_L_0_out, I1 =>  C_48_S_0_L_1_out, I2 =>  C_48_S_0_L_2_out, I3 =>  C_48_S_0_L_3_out, I4 =>  C_48_S_0_L_4_out, I5 =>  C_48_S_0_L_5_out, I6 =>  C_48_S_0_L_6_out, I7 =>  C_48_S_0_L_7_out); 
C_48_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111111101110100011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100011101000100000001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_48_S_1_out, I0 =>  C_48_S_1_L_0_out, I1 =>  C_48_S_1_L_1_out, I2 =>  C_48_S_1_L_2_out, I3 =>  C_48_S_1_L_3_out, I4 =>  C_48_S_1_L_4_out, I5 =>  C_48_S_1_L_5_out, I6 =>  C_48_S_1_L_6_out, I7 =>  C_48_S_1_L_7_out); 
C_48_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110101010101000111111101110101011101010101010001110101010101000111010001000000011111110111010001110101010101000111010101010100010101000100000001110101010101000111010001000000011101000100000001000000000000000") port map( O =>C_48_S_2_out, I0 =>  C_48_S_2_L_0_out, I1 =>  C_48_S_2_L_1_out, I2 =>  C_48_S_2_L_2_out, I3 =>  C_48_S_2_L_3_out, I4 =>  C_48_S_2_L_4_out, I5 =>  C_48_S_2_L_5_out, I6 =>  C_48_S_2_L_6_out, I7 =>  C_48_S_2_L_7_out); 
C_48_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111111101110101011101010101010001110101010001000101010001000000011111110111010101110111010101000111010101010100010101000100000001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_48_S_3_out, I0 =>  C_48_S_3_L_0_out, I1 =>  C_48_S_3_L_1_out, I2 =>  C_48_S_3_L_2_out, I3 =>  C_48_S_3_L_3_out, I4 =>  C_48_S_3_L_4_out, I5 =>  C_48_S_3_L_5_out, I6 =>  C_48_S_3_L_6_out, I7 =>  C_48_S_3_L_7_out); 
C_48_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101111110011111110111111001111110011001000111111101111110011111100110000001111110011101000110000001000000011111110111111001110100011000000111111001100000011000000100000001110110011000000110000001000000011000000100000001000000000000000") port map( O =>C_48_S_4_out, I0 =>  C_48_S_4_L_0_out, I1 =>  C_48_S_4_L_1_out, I2 =>  C_48_S_4_L_2_out, I3 =>  C_48_S_4_L_3_out, I4 =>  C_48_S_4_L_4_out, I5 =>  C_48_S_4_L_5_out, I6 =>  C_48_S_4_L_6_out, I7 =>  C_48_S_4_L_7_out); 

C_48_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_48_out, I0 =>  C_48_S_0_out, I1 =>  C_48_S_1_out, I2 =>  C_48_S_2_out, I3 =>  C_48_S_3_out, I4 =>  C_48_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_49_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101110101011101010101010101110101010101010111010101010101010101010101010001010101010101000101010001010100011101010111010101110101010101010111010101010101010101010101010001010101010101000101010101010100010101000101010001010100010001000") port map( O =>C_49_S_0_out, I0 =>  C_49_S_0_L_0_out, I1 =>  C_49_S_0_L_1_out, I2 =>  C_49_S_0_L_2_out, I3 =>  C_49_S_0_L_3_out, I4 =>  C_49_S_0_L_4_out, I5 =>  C_49_S_0_L_5_out, I6 =>  C_49_S_0_L_6_out, I7 =>  C_49_S_0_L_7_out); 
C_49_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010001110101011101000111111101110101011101010111010001110101011101000111010001000000011111110111010001110100010101000111010001010100010101000100000001110100010101000111010001000000010101000100000001000000000000000") port map( O =>C_49_S_1_out, I0 =>  C_49_S_1_L_0_out, I1 =>  C_49_S_1_L_1_out, I2 =>  C_49_S_1_L_2_out, I3 =>  C_49_S_1_L_3_out, I4 =>  C_49_S_1_L_4_out, I5 =>  C_49_S_1_L_5_out, I6 =>  C_49_S_1_L_6_out, I7 =>  C_49_S_1_L_7_out); 
C_49_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001111110011001000111111101110100011111110111010001110100011000000111010001000000011111110111010001111110011101000111010001000000011101000100000001110110011000000111010001000000011101000100000001000000000000000") port map( O =>C_49_S_2_out, I0 =>  C_49_S_2_L_0_out, I1 =>  C_49_S_2_L_1_out, I2 =>  C_49_S_2_L_2_out, I3 =>  C_49_S_2_L_3_out, I4 =>  C_49_S_2_L_4_out, I5 =>  C_49_S_2_L_5_out, I6 =>  C_49_S_2_L_6_out, I7 =>  C_49_S_2_L_7_out); 
C_49_S_3_inst : LUT8 generic map(INIT => "1111111111101110111011101110100011111110111010001110100010001000111111101110110011101100100010001110111011001000110010001000000011111110111011001110110010001000111011101100100011001000100000001110111011101000111010001000000011101000100010001000100000000000") port map( O =>C_49_S_3_out, I0 =>  C_49_S_3_L_0_out, I1 =>  C_49_S_3_L_1_out, I2 =>  C_49_S_3_L_2_out, I3 =>  C_49_S_3_L_3_out, I4 =>  C_49_S_3_L_4_out, I5 =>  C_49_S_3_L_5_out, I6 =>  C_49_S_3_L_6_out, I7 =>  C_49_S_3_L_7_out); 
C_49_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_49_S_4_out, I0 =>  C_49_S_4_L_0_out, I1 =>  C_49_S_4_L_1_out, I2 =>  C_49_S_4_L_2_out, I3 =>  C_49_S_4_L_3_out, I4 =>  C_49_S_4_L_4_out, I5 =>  C_49_S_4_L_5_out, I6 =>  C_49_S_4_L_6_out, I7 =>  C_49_S_4_L_7_out); 

C_49_inst : LUT8 generic map(INIT => "1110101011101010101010001010100011101010111010101010100010101000111010101110101010101000101010001110101011101010101010001010100011101010111010101010100010101000111010101110101010101000101010001110101011101010101010001010100011101010111010101010100010101000") port map( O =>C_49_out, I0 =>  C_49_S_0_out, I1 =>  C_49_S_1_out, I2 =>  C_49_S_2_out, I3 =>  C_49_S_3_out, I4 =>  C_49_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_50_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101010111010101110101010101010111010101010101010101010101010001010101010101010101010001010100011101010111010101010101010101010111010101010101010101010101010001010101010101000101010001010100010101010101010001010100010001000") port map( O =>C_50_S_0_out, I0 =>  C_50_S_0_L_0_out, I1 =>  C_50_S_0_L_1_out, I2 =>  C_50_S_0_L_2_out, I3 =>  C_50_S_0_L_3_out, I4 =>  C_50_S_0_L_4_out, I5 =>  C_50_S_0_L_5_out, I6 =>  C_50_S_0_L_6_out, I7 =>  C_50_S_0_L_7_out); 
C_50_S_1_inst : LUT8 generic map(INIT => "1111111111101110111011101010101011111110111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001000000010101010100010001000100000000000") port map( O =>C_50_S_1_out, I0 =>  C_50_S_1_L_0_out, I1 =>  C_50_S_1_L_1_out, I2 =>  C_50_S_1_L_2_out, I3 =>  C_50_S_1_L_3_out, I4 =>  C_50_S_1_L_4_out, I5 =>  C_50_S_1_L_5_out, I6 =>  C_50_S_1_L_6_out, I7 =>  C_50_S_1_L_7_out); 
C_50_S_2_inst : LUT8 generic map(INIT => "1111111111111110111110101110100011111110111110101110100010100000111110101111101010101000101000001110100010101000100000001000000011111110111111101110101011101000111110101110101010100000101000001111101011101000101000001000000011101000101000001000000000000000") port map( O =>C_50_S_2_out, I0 =>  C_50_S_2_L_0_out, I1 =>  C_50_S_2_L_1_out, I2 =>  C_50_S_2_L_2_out, I3 =>  C_50_S_2_L_3_out, I4 =>  C_50_S_2_L_4_out, I5 =>  C_50_S_2_L_5_out, I6 =>  C_50_S_2_L_6_out, I7 =>  C_50_S_2_L_7_out); 
C_50_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111110111011111111111111101110111010001000111111111111111011101100100000001111111011101000100000000000000011111111111111101110100010000000111111101100100010000000000000001110111010001000100000000000000010001000000000000000000000000000") port map( O =>C_50_S_3_out, I0 =>  C_50_S_3_L_0_out, I1 =>  C_50_S_3_L_1_out, I2 =>  C_50_S_3_L_2_out, I3 =>  C_50_S_3_L_3_out, I4 =>  C_50_S_3_L_4_out, I5 =>  C_50_S_3_L_5_out, I6 =>  C_50_S_3_L_6_out, I7 =>  C_50_S_3_L_7_out); 
C_50_S_4_inst : LUT8 generic map(INIT => "1111111011111100111111101110100011111110111010001111100011100000111111101110100011111000111010001111111011101000111010001000000011111110111010001110100010000000111010001110000011101000100000001111100011100000111010001000000011101000100000001100000010000000") port map( O =>C_50_S_4_out, I0 =>  C_50_S_4_L_0_out, I1 =>  C_50_S_4_L_1_out, I2 =>  C_50_S_4_L_2_out, I3 =>  C_50_S_4_L_3_out, I4 =>  C_50_S_4_L_4_out, I5 =>  C_50_S_4_L_5_out, I6 =>  C_50_S_4_L_6_out, I7 =>  C_50_S_4_L_7_out); 

C_50_inst : LUT8 generic map(INIT => "1110101010101010101010101010100011101010101010101010101010101000111010101010101010101010101010001110101010101010101010101010100011101010101010101010101010101000111010101010101010101010101010001110101010101010101010101010100011101010101010101010101010101000") port map( O =>C_50_out, I0 =>  C_50_S_0_out, I1 =>  C_50_S_1_out, I2 =>  C_50_S_2_out, I3 =>  C_50_S_3_out, I4 =>  C_50_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_51_S_0_inst : LUT8 generic map(INIT => "1110111011101010111011101110101011101010111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001010100010101000100010001010100010001000") port map( O =>C_51_S_0_out, I0 =>  C_51_S_0_L_0_out, I1 =>  C_51_S_0_L_1_out, I2 =>  C_51_S_0_L_2_out, I3 =>  C_51_S_0_L_3_out, I4 =>  C_51_S_0_L_4_out, I5 =>  C_51_S_0_L_5_out, I6 =>  C_51_S_0_L_6_out, I7 =>  C_51_S_0_L_7_out); 
C_51_S_1_inst : LUT8 generic map(INIT => "1111111011111010111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001010000011111010111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001010000010000000") port map( O =>C_51_S_1_out, I0 =>  C_51_S_1_L_0_out, I1 =>  C_51_S_1_L_1_out, I2 =>  C_51_S_1_L_2_out, I3 =>  C_51_S_1_L_3_out, I4 =>  C_51_S_1_L_4_out, I5 =>  C_51_S_1_L_5_out, I6 =>  C_51_S_1_L_6_out, I7 =>  C_51_S_1_L_7_out); 
C_51_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110110011111110111010001110100011001000111111101111111011101110111010001110100011101000111010001000000011111110111010001110100011101000111010001000100010000000100000001110110011101000111010001000000011001000100000001000000000000000") port map( O =>C_51_S_2_out, I0 =>  C_51_S_2_L_0_out, I1 =>  C_51_S_2_L_1_out, I2 =>  C_51_S_2_L_2_out, I3 =>  C_51_S_2_L_3_out, I4 =>  C_51_S_2_L_4_out, I5 =>  C_51_S_2_L_5_out, I6 =>  C_51_S_2_L_6_out, I7 =>  C_51_S_2_L_7_out); 
C_51_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_51_S_3_out, I0 =>  C_51_S_3_L_0_out, I1 =>  C_51_S_3_L_1_out, I2 =>  C_51_S_3_L_2_out, I3 =>  C_51_S_3_L_3_out, I4 =>  C_51_S_3_L_4_out, I5 =>  C_51_S_3_L_5_out, I6 =>  C_51_S_3_L_6_out, I7 =>  C_51_S_3_L_7_out); 
C_51_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111101110111011111110111010001110111010101000111010001000000011111110111010001110101010001000111010001000000010001000100000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_51_S_4_out, I0 =>  C_51_S_4_L_0_out, I1 =>  C_51_S_4_L_1_out, I2 =>  C_51_S_4_L_2_out, I3 =>  C_51_S_4_L_3_out, I4 =>  C_51_S_4_L_4_out, I5 =>  C_51_S_4_L_5_out, I6 =>  C_51_S_4_L_6_out, I7 =>  C_51_S_4_L_7_out); 

C_51_inst : LUT8 generic map(INIT => "1110101011101010101010001010100011101010111010101010100010101000111010101110101010101000101010001110101011101010101010001010100011101010111010101010100010101000111010101110101010101000101010001110101011101010101010001010100011101010111010101010100010101000") port map( O =>C_51_out, I0 =>  C_51_S_0_out, I1 =>  C_51_S_1_out, I2 =>  C_51_S_2_out, I3 =>  C_51_S_3_out, I4 =>  C_51_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_52_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010100011101010101010101010101010101010101010101010101010101010101010001010101010101010101010101010100010101010101010001010100010001000") port map( O =>C_52_S_0_out, I0 =>  C_52_S_0_L_0_out, I1 =>  C_52_S_0_L_1_out, I2 =>  C_52_S_0_L_2_out, I3 =>  C_52_S_0_L_3_out, I4 =>  C_52_S_0_L_4_out, I5 =>  C_52_S_0_L_5_out, I6 =>  C_52_S_0_L_6_out, I7 =>  C_52_S_0_L_7_out); 
C_52_S_1_inst : LUT8 generic map(INIT => "1111111011101110111111101110101011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100010101000100000001000100010000000") port map( O =>C_52_S_1_out, I0 =>  C_52_S_1_L_0_out, I1 =>  C_52_S_1_L_1_out, I2 =>  C_52_S_1_L_2_out, I3 =>  C_52_S_1_L_3_out, I4 =>  C_52_S_1_L_4_out, I5 =>  C_52_S_1_L_5_out, I6 =>  C_52_S_1_L_6_out, I7 =>  C_52_S_1_L_7_out); 
C_52_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111011101110111011101000111111101110110011101100111010001110100011101000110010001000000011111110111011001110100011101000111010001100100011001000100000001110100010001000100010001000000010001000100000001000000000000000") port map( O =>C_52_S_2_out, I0 =>  C_52_S_2_L_0_out, I1 =>  C_52_S_2_L_1_out, I2 =>  C_52_S_2_L_2_out, I3 =>  C_52_S_2_L_3_out, I4 =>  C_52_S_2_L_4_out, I5 =>  C_52_S_2_L_5_out, I6 =>  C_52_S_2_L_6_out, I7 =>  C_52_S_2_L_7_out); 
C_52_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111110111111001111110011101000111111101111110011111100111010001111100011000000110000001000000011111110111111001111110011100000111010001100000011000000100000001110100011000000110000001000000011000000000000000000000000000000") port map( O =>C_52_S_3_out, I0 =>  C_52_S_3_L_0_out, I1 =>  C_52_S_3_L_1_out, I2 =>  C_52_S_3_L_2_out, I3 =>  C_52_S_3_L_3_out, I4 =>  C_52_S_3_L_4_out, I5 =>  C_52_S_3_L_5_out, I6 =>  C_52_S_3_L_6_out, I7 =>  C_52_S_3_L_7_out); 
C_52_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101111110011111110111111001111110011101000111111101111110011111000110000001111110011100000110000001000000011111110111111001111100011000000111111001110000011000000100000001110100011000000110000001000000011000000100000001000000000000000") port map( O =>C_52_S_4_out, I0 =>  C_52_S_4_L_0_out, I1 =>  C_52_S_4_L_1_out, I2 =>  C_52_S_4_L_2_out, I3 =>  C_52_S_4_L_3_out, I4 =>  C_52_S_4_L_4_out, I5 =>  C_52_S_4_L_5_out, I6 =>  C_52_S_4_L_6_out, I7 =>  C_52_S_4_L_7_out); 

C_52_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_52_out, I0 =>  C_52_S_0_out, I1 =>  C_52_S_1_out, I2 =>  C_52_S_2_out, I3 =>  C_52_S_3_out, I4 =>  C_52_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_53_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_53_S_0_out, I0 =>  C_53_S_0_L_0_out, I1 =>  C_53_S_0_L_1_out, I2 =>  C_53_S_0_L_2_out, I3 =>  C_53_S_0_L_3_out, I4 =>  C_53_S_0_L_4_out, I5 =>  C_53_S_0_L_5_out, I6 =>  C_53_S_0_L_6_out, I7 =>  C_53_S_0_L_7_out); 
C_53_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_53_S_1_out, I0 =>  C_53_S_1_L_0_out, I1 =>  C_53_S_1_L_1_out, I2 =>  C_53_S_1_L_2_out, I3 =>  C_53_S_1_L_3_out, I4 =>  C_53_S_1_L_4_out, I5 =>  C_53_S_1_L_5_out, I6 =>  C_53_S_1_L_6_out, I7 =>  C_53_S_1_L_7_out); 
C_53_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_53_S_2_out, I0 =>  C_53_S_2_L_0_out, I1 =>  C_53_S_2_L_1_out, I2 =>  C_53_S_2_L_2_out, I3 =>  C_53_S_2_L_3_out, I4 =>  C_53_S_2_L_4_out, I5 =>  C_53_S_2_L_5_out, I6 =>  C_53_S_2_L_6_out, I7 =>  C_53_S_2_L_7_out); 
C_53_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_53_S_3_out, I0 =>  C_53_S_3_L_0_out, I1 =>  C_53_S_3_L_1_out, I2 =>  C_53_S_3_L_2_out, I3 =>  C_53_S_3_L_3_out, I4 =>  C_53_S_3_L_4_out, I5 =>  C_53_S_3_L_5_out, I6 =>  C_53_S_3_L_6_out, I7 =>  C_53_S_3_L_7_out); 
C_53_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_53_S_4_out, I0 =>  C_53_S_4_L_0_out, I1 =>  C_53_S_4_L_1_out, I2 =>  C_53_S_4_L_2_out, I3 =>  C_53_S_4_L_3_out, I4 =>  C_53_S_4_L_4_out, I5 =>  C_53_S_4_L_5_out, I6 =>  C_53_S_4_L_6_out, I7 =>  C_53_S_4_L_7_out); 

C_53_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_53_out, I0 =>  C_53_S_0_out, I1 =>  C_53_S_1_out, I2 =>  C_53_S_2_out, I3 =>  C_53_S_3_out, I4 =>  C_53_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_54_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101010101010101010101010101000111010101010101011101010101010101010101010101000101010101010100011101010101010101110101010101010101010101010100010101010101010001110101010101010101010101010100010101010101010001010100010001000") port map( O =>C_54_S_0_out, I0 =>  C_54_S_0_L_0_out, I1 =>  C_54_S_0_L_1_out, I2 =>  C_54_S_0_L_2_out, I3 =>  C_54_S_0_L_3_out, I4 =>  C_54_S_0_L_4_out, I5 =>  C_54_S_0_L_5_out, I6 =>  C_54_S_0_L_6_out, I7 =>  C_54_S_0_L_7_out); 
C_54_S_1_inst : LUT8 generic map(INIT => "1111111011111010111111101110101011111010111010101110101010101000111110101110100011101010101010001110100010101000101010001000000011111110111010101110101011101000111010101010100011101000101000001110101010101000101010001010000010101000100000001010000010000000") port map( O =>C_54_S_1_out, I0 =>  C_54_S_1_L_0_out, I1 =>  C_54_S_1_L_1_out, I2 =>  C_54_S_1_L_2_out, I3 =>  C_54_S_1_L_3_out, I4 =>  C_54_S_1_L_4_out, I5 =>  C_54_S_1_L_5_out, I6 =>  C_54_S_1_L_6_out, I7 =>  C_54_S_1_L_7_out); 
C_54_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010100000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001111101011101000111010001000000011101000100000001000000000000000") port map( O =>C_54_S_2_out, I0 =>  C_54_S_2_L_0_out, I1 =>  C_54_S_2_L_1_out, I2 =>  C_54_S_2_L_2_out, I3 =>  C_54_S_2_L_3_out, I4 =>  C_54_S_2_L_4_out, I5 =>  C_54_S_2_L_5_out, I6 =>  C_54_S_2_L_6_out, I7 =>  C_54_S_2_L_7_out); 
C_54_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010100000101000001000000011111110111110101111101011101000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_54_S_3_out, I0 =>  C_54_S_3_L_0_out, I1 =>  C_54_S_3_L_1_out, I2 =>  C_54_S_3_L_2_out, I3 =>  C_54_S_3_L_3_out, I4 =>  C_54_S_3_L_4_out, I5 =>  C_54_S_3_L_5_out, I6 =>  C_54_S_3_L_6_out, I7 =>  C_54_S_3_L_7_out); 
C_54_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101111111011111110111111101110111011101000111111101110110011101000110010001110100011001000110010001000000011111110111011001110110011101000111011001110100011001000100000001110100010001000100000001000000010000000100000001000000000000000") port map( O =>C_54_S_4_out, I0 =>  C_54_S_4_L_0_out, I1 =>  C_54_S_4_L_1_out, I2 =>  C_54_S_4_L_2_out, I3 =>  C_54_S_4_L_3_out, I4 =>  C_54_S_4_L_4_out, I5 =>  C_54_S_4_L_5_out, I6 =>  C_54_S_4_L_6_out, I7 =>  C_54_S_4_L_7_out); 

C_54_inst : LUT8 generic map(INIT => "1110101011101000111010001010100011101010111010001110100010101000111010101110100011101000101010001110101011101000111010001010100011101010111010001110100010101000111010101110100011101000101010001110101011101000111010001010100011101010111010001110100010101000") port map( O =>C_54_out, I0 =>  C_54_S_0_out, I1 =>  C_54_S_1_out, I2 =>  C_54_S_2_out, I3 =>  C_54_S_3_out, I4 =>  C_54_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_55_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101010101010101010101010101000111010101010101010101010101010001110101010101010101010101010100011101010101010101010101010101000111010101010101010101010101010001110101010101010101010101010100010101010101010001010100010001000") port map( O =>C_55_S_0_out, I0 =>  C_55_S_0_L_0_out, I1 =>  C_55_S_0_L_1_out, I2 =>  C_55_S_0_L_2_out, I3 =>  C_55_S_0_L_3_out, I4 =>  C_55_S_0_L_4_out, I5 =>  C_55_S_0_L_5_out, I6 =>  C_55_S_0_L_6_out, I7 =>  C_55_S_0_L_7_out); 
C_55_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010101110101010101000111111101110101011101010101010001110111010101000101010001000000011111110111010101110101010001000111010101010100010101000100000001110101010101000101010001000000011101000100000001000000000000000") port map( O =>C_55_S_1_out, I0 =>  C_55_S_1_L_0_out, I1 =>  C_55_S_1_L_1_out, I2 =>  C_55_S_1_L_2_out, I3 =>  C_55_S_1_L_3_out, I4 =>  C_55_S_1_L_4_out, I5 =>  C_55_S_1_L_5_out, I6 =>  C_55_S_1_L_6_out, I7 =>  C_55_S_1_L_7_out); 
C_55_S_2_inst : LUT8 generic map(INIT => "1111111111111100111111101110100011111110111010001111110011000000111111101110100011111100110000001111110011000000111010001000000011111110111010001111110011000000111111001100000011101000100000001111110011000000111010001000000011101000100000001100000000000000") port map( O =>C_55_S_2_out, I0 =>  C_55_S_2_L_0_out, I1 =>  C_55_S_2_L_1_out, I2 =>  C_55_S_2_L_2_out, I3 =>  C_55_S_2_L_3_out, I4 =>  C_55_S_2_L_4_out, I5 =>  C_55_S_2_L_5_out, I6 =>  C_55_S_2_L_6_out, I7 =>  C_55_S_2_L_7_out); 
C_55_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111110101110100010100000111111111111111011111010111010001111111011101000111010001000000011111110111010001110100010000000111010001010000010000000000000001111101011101000101000001000000011101000100000001000000000000000") port map( O =>C_55_S_3_out, I0 =>  C_55_S_3_L_0_out, I1 =>  C_55_S_3_L_1_out, I2 =>  C_55_S_3_L_2_out, I3 =>  C_55_S_3_L_3_out, I4 =>  C_55_S_3_L_4_out, I5 =>  C_55_S_3_L_5_out, I6 =>  C_55_S_3_L_6_out, I7 =>  C_55_S_3_L_7_out); 
C_55_S_4_inst : LUT8 generic map(INIT => "1111111111111010111111101110100011111110111010001110100010100000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001111101011101000111010001000000011101000100000001010000000000000") port map( O =>C_55_S_4_out, I0 =>  C_55_S_4_L_0_out, I1 =>  C_55_S_4_L_1_out, I2 =>  C_55_S_4_L_2_out, I3 =>  C_55_S_4_L_3_out, I4 =>  C_55_S_4_L_4_out, I5 =>  C_55_S_4_L_5_out, I6 =>  C_55_S_4_L_6_out, I7 =>  C_55_S_4_L_7_out); 

C_55_inst : LUT8 generic map(INIT => "1110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000") port map( O =>C_55_out, I0 =>  C_55_S_0_out, I1 =>  C_55_S_1_out, I2 =>  C_55_S_2_out, I3 =>  C_55_S_3_out, I4 =>  C_55_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_56_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111000111000001111100010100000100000000000000011111111111111101111101011100000111110001110000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_56_S_0_out, I0 =>  C_56_S_0_L_0_out, I1 =>  C_56_S_0_L_1_out, I2 =>  C_56_S_0_L_2_out, I3 =>  C_56_S_0_L_3_out, I4 =>  C_56_S_0_L_4_out, I5 =>  C_56_S_0_L_5_out, I6 =>  C_56_S_0_L_6_out, I7 =>  C_56_S_0_L_7_out); 
C_56_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111110111010001111111011100000111000001000000011111110111110001111100010000000111010001000000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_56_S_1_out, I0 =>  C_56_S_1_L_0_out, I1 =>  C_56_S_1_L_1_out, I2 =>  C_56_S_1_L_2_out, I3 =>  C_56_S_1_L_3_out, I4 =>  C_56_S_1_L_4_out, I5 =>  C_56_S_1_L_5_out, I6 =>  C_56_S_1_L_6_out, I7 =>  C_56_S_1_L_7_out); 
C_56_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_56_S_2_out, I0 =>  C_56_S_2_L_0_out, I1 =>  C_56_S_2_L_1_out, I2 =>  C_56_S_2_L_2_out, I3 =>  C_56_S_2_L_3_out, I4 =>  C_56_S_2_L_4_out, I5 =>  C_56_S_2_L_5_out, I6 =>  C_56_S_2_L_6_out, I7 =>  C_56_S_2_L_7_out); 
C_56_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111100010000000100000000000000011111111111111101111111011100000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_56_S_3_out, I0 =>  C_56_S_3_L_0_out, I1 =>  C_56_S_3_L_1_out, I2 =>  C_56_S_3_L_2_out, I3 =>  C_56_S_3_L_3_out, I4 =>  C_56_S_3_L_4_out, I5 =>  C_56_S_3_L_5_out, I6 =>  C_56_S_3_L_6_out, I7 =>  C_56_S_3_L_7_out); 
C_56_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_56_S_4_out, I0 =>  C_56_S_4_L_0_out, I1 =>  C_56_S_4_L_1_out, I2 =>  C_56_S_4_L_2_out, I3 =>  C_56_S_4_L_3_out, I4 =>  C_56_S_4_L_4_out, I5 =>  C_56_S_4_L_5_out, I6 =>  C_56_S_4_L_6_out, I7 =>  C_56_S_4_L_7_out); 

C_56_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_56_out, I0 =>  C_56_S_0_out, I1 =>  C_56_S_1_out, I2 =>  C_56_S_2_out, I3 =>  C_56_S_3_out, I4 =>  C_56_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_57_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_57_S_0_out, I0 =>  C_57_S_0_L_0_out, I1 =>  C_57_S_0_L_1_out, I2 =>  C_57_S_0_L_2_out, I3 =>  C_57_S_0_L_3_out, I4 =>  C_57_S_0_L_4_out, I5 =>  C_57_S_0_L_5_out, I6 =>  C_57_S_0_L_6_out, I7 =>  C_57_S_0_L_7_out); 
C_57_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_57_S_1_out, I0 =>  C_57_S_1_L_0_out, I1 =>  C_57_S_1_L_1_out, I2 =>  C_57_S_1_L_2_out, I3 =>  C_57_S_1_L_3_out, I4 =>  C_57_S_1_L_4_out, I5 =>  C_57_S_1_L_5_out, I6 =>  C_57_S_1_L_6_out, I7 =>  C_57_S_1_L_7_out); 
C_57_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_57_S_2_out, I0 =>  C_57_S_2_L_0_out, I1 =>  C_57_S_2_L_1_out, I2 =>  C_57_S_2_L_2_out, I3 =>  C_57_S_2_L_3_out, I4 =>  C_57_S_2_L_4_out, I5 =>  C_57_S_2_L_5_out, I6 =>  C_57_S_2_L_6_out, I7 =>  C_57_S_2_L_7_out); 
C_57_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_57_S_3_out, I0 =>  C_57_S_3_L_0_out, I1 =>  C_57_S_3_L_1_out, I2 =>  C_57_S_3_L_2_out, I3 =>  C_57_S_3_L_3_out, I4 =>  C_57_S_3_L_4_out, I5 =>  C_57_S_3_L_5_out, I6 =>  C_57_S_3_L_6_out, I7 =>  C_57_S_3_L_7_out); 
C_57_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111110011111111111111001111110011000000111111111111110011111100110000001111110011000000110000000000000011111111111111001111110011000000111111001100000011000000000000001111110011000000110000000000000011000000000000000000000000000000") port map( O =>C_57_S_4_out, I0 =>  C_57_S_4_L_0_out, I1 =>  C_57_S_4_L_1_out, I2 =>  C_57_S_4_L_2_out, I3 =>  C_57_S_4_L_3_out, I4 =>  C_57_S_4_L_4_out, I5 =>  C_57_S_4_L_5_out, I6 =>  C_57_S_4_L_6_out, I7 =>  C_57_S_4_L_7_out); 

C_57_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_57_out, I0 =>  C_57_S_0_out, I1 =>  C_57_S_1_out, I2 =>  C_57_S_2_out, I3 =>  C_57_S_3_out, I4 =>  C_57_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_58_S_0_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110101011101000111111101110100011101000101000001110100010101000111010001000000011111110111010001110101011101000111110101110100011101000100000001110100010101000111010001000000011101000100000001000000010000000") port map( O =>C_58_S_0_out, I0 =>  C_58_S_0_L_0_out, I1 =>  C_58_S_0_L_1_out, I2 =>  C_58_S_0_L_2_out, I3 =>  C_58_S_0_L_3_out, I4 =>  C_58_S_0_L_4_out, I5 =>  C_58_S_0_L_5_out, I6 =>  C_58_S_0_L_6_out, I7 =>  C_58_S_0_L_7_out); 
C_58_S_1_inst : LUT8 generic map(INIT => "1111111111101010111111101110100011111110111010001111101010101000111111101110100011101010101000001111101010101000111010001000000011111110111010001110101010100000111110101010100011101000100000001110101010100000111010001000000011101000100000001010100000000000") port map( O =>C_58_S_1_out, I0 =>  C_58_S_1_L_0_out, I1 =>  C_58_S_1_L_1_out, I2 =>  C_58_S_1_L_2_out, I3 =>  C_58_S_1_L_3_out, I4 =>  C_58_S_1_L_4_out, I5 =>  C_58_S_1_L_5_out, I6 =>  C_58_S_1_L_6_out, I7 =>  C_58_S_1_L_7_out); 
C_58_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110111010001000111111101110101011101010100010001110111010001000101010000000000011111111111010101110111010001000111011101010100010101000100000001110111010001000101010001000000010101000100000001000000000000000") port map( O =>C_58_S_2_out, I0 =>  C_58_S_2_L_0_out, I1 =>  C_58_S_2_L_1_out, I2 =>  C_58_S_2_L_2_out, I3 =>  C_58_S_2_L_3_out, I4 =>  C_58_S_2_L_4_out, I5 =>  C_58_S_2_L_5_out, I6 =>  C_58_S_2_L_6_out, I7 =>  C_58_S_2_L_7_out); 
C_58_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010101110100011101000111111101110101011101000111010001111101011101000111010001000000011111110111010001110100010100000111010001110100010101000100000001110100011101000101010001000000011101000100000001000000000000000") port map( O =>C_58_S_3_out, I0 =>  C_58_S_3_L_0_out, I1 =>  C_58_S_3_L_1_out, I2 =>  C_58_S_3_L_2_out, I3 =>  C_58_S_3_L_3_out, I4 =>  C_58_S_3_L_4_out, I5 =>  C_58_S_3_L_5_out, I6 =>  C_58_S_3_L_6_out, I7 =>  C_58_S_3_L_7_out); 
C_58_S_4_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110101011101000111010001000000011111110111010001110100010101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_58_S_4_out, I0 =>  C_58_S_4_L_0_out, I1 =>  C_58_S_4_L_1_out, I2 =>  C_58_S_4_L_2_out, I3 =>  C_58_S_4_L_3_out, I4 =>  C_58_S_4_L_4_out, I5 =>  C_58_S_4_L_5_out, I6 =>  C_58_S_4_L_6_out, I7 =>  C_58_S_4_L_7_out); 

C_58_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_58_out, I0 =>  C_58_S_0_out, I1 =>  C_58_S_1_out, I2 =>  C_58_S_2_out, I3 =>  C_58_S_3_out, I4 =>  C_58_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_59_S_0_inst : LUT8 generic map(INIT => "1110111011101010111010101010101011101010101010101110101010101000111010101010101011101010101010001110101010101000101010101010100011101010101010101110101010101000111010101010100010101010101010001110101010101000101010101010100010101010101010001010100010001000") port map( O =>C_59_S_0_out, I0 =>  C_59_S_0_L_0_out, I1 =>  C_59_S_0_L_1_out, I2 =>  C_59_S_0_L_2_out, I3 =>  C_59_S_0_L_3_out, I4 =>  C_59_S_0_L_4_out, I5 =>  C_59_S_0_L_5_out, I6 =>  C_59_S_0_L_6_out, I7 =>  C_59_S_0_L_7_out); 
C_59_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101110100011111110111010101110100010101000111111101110100011101000101010001110101011101000101010001000000011111110111010101110100010101000111010101110100011101000100000001110101011101000101010001000000011101000101010001010100010000000") port map( O =>C_59_S_1_out, I0 =>  C_59_S_1_L_0_out, I1 =>  C_59_S_1_L_1_out, I2 =>  C_59_S_1_L_2_out, I3 =>  C_59_S_1_L_3_out, I4 =>  C_59_S_1_L_4_out, I5 =>  C_59_S_1_L_5_out, I6 =>  C_59_S_1_L_6_out, I7 =>  C_59_S_1_L_7_out); 
C_59_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111011101110111011101000111111101110110011101100111010001110110011101000111010001000000011111110111010001110100011001000111010001100100011001000100000001110100010001000100010001000000010001000100000001000000000000000") port map( O =>C_59_S_2_out, I0 =>  C_59_S_2_L_0_out, I1 =>  C_59_S_2_L_1_out, I2 =>  C_59_S_2_L_2_out, I3 =>  C_59_S_2_L_3_out, I4 =>  C_59_S_2_L_4_out, I5 =>  C_59_S_2_L_5_out, I6 =>  C_59_S_2_L_6_out, I7 =>  C_59_S_2_L_7_out); 
C_59_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111111111110011111111111011001111110011000000111111101110100011111100110000001111110011000000111010001000000011111110111010001111110011000000111111001100000011101000100000001111110011000000110010000000000011000000000000001000000000000000") port map( O =>C_59_S_3_out, I0 =>  C_59_S_3_L_0_out, I1 =>  C_59_S_3_L_1_out, I2 =>  C_59_S_3_L_2_out, I3 =>  C_59_S_3_L_3_out, I4 =>  C_59_S_3_L_4_out, I5 =>  C_59_S_3_L_5_out, I6 =>  C_59_S_3_L_6_out, I7 =>  C_59_S_3_L_7_out); 
C_59_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111111110111011111110111010101111111011101000111111101110100011101010100010001110101010000000101010001000000011111110111010101111111010101000111011101010100011101000100000001110100010000000101010001000000010001000000000001000000000000000") port map( O =>C_59_S_4_out, I0 =>  C_59_S_4_L_0_out, I1 =>  C_59_S_4_L_1_out, I2 =>  C_59_S_4_L_2_out, I3 =>  C_59_S_4_L_3_out, I4 =>  C_59_S_4_L_4_out, I5 =>  C_59_S_4_L_5_out, I6 =>  C_59_S_4_L_6_out, I7 =>  C_59_S_4_L_7_out); 

C_59_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_59_out, I0 =>  C_59_S_0_out, I1 =>  C_59_S_1_out, I2 =>  C_59_S_2_out, I3 =>  C_59_S_3_out, I4 =>  C_59_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_60_S_0_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_60_S_0_out, I0 =>  C_60_S_0_L_0_out, I1 =>  C_60_S_0_L_1_out, I2 =>  C_60_S_0_L_2_out, I3 =>  C_60_S_0_L_3_out, I4 =>  C_60_S_0_L_4_out, I5 =>  C_60_S_0_L_5_out, I6 =>  C_60_S_0_L_6_out, I7 =>  C_60_S_0_L_7_out); 
C_60_S_1_inst : LUT8 generic map(INIT => "1111111011101000111111101110100011111110111010001111111010000000111111101110100011111110100000001111101010000000111010001000000011111110111010001111111010100000111111101000000011101000100000001111111010000000111010001000000011101000100000001110100010000000") port map( O =>C_60_S_1_out, I0 =>  C_60_S_1_L_0_out, I1 =>  C_60_S_1_L_1_out, I2 =>  C_60_S_1_L_2_out, I3 =>  C_60_S_1_L_3_out, I4 =>  C_60_S_1_L_4_out, I5 =>  C_60_S_1_L_5_out, I6 =>  C_60_S_1_L_6_out, I7 =>  C_60_S_1_L_7_out); 
C_60_S_2_inst : LUT8 generic map(INIT => "1111111011101000111111101110100011111110111010001110100010000000111111101110100011111110111010001111101010000000111010001000000011111110111010001111111010100000111010001000000011101000100000001111111011101000111010001000000011101000100000001110100010000000") port map( O =>C_60_S_2_out, I0 =>  C_60_S_2_L_0_out, I1 =>  C_60_S_2_L_1_out, I2 =>  C_60_S_2_L_2_out, I3 =>  C_60_S_2_L_3_out, I4 =>  C_60_S_2_L_4_out, I5 =>  C_60_S_2_L_5_out, I6 =>  C_60_S_2_L_6_out, I7 =>  C_60_S_2_L_7_out); 
C_60_S_3_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110111011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100010001000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_60_S_3_out, I0 =>  C_60_S_3_L_0_out, I1 =>  C_60_S_3_L_1_out, I2 =>  C_60_S_3_L_2_out, I3 =>  C_60_S_3_L_3_out, I4 =>  C_60_S_3_L_4_out, I5 =>  C_60_S_3_L_5_out, I6 =>  C_60_S_3_L_6_out, I7 =>  C_60_S_3_L_7_out); 
C_60_S_4_inst : LUT8 generic map(INIT => "1111111011101000111111101110100011111110111010001111111011101000111111101110100011111010111010001111101011101000111010001000000011111110111010001110100010100000111010001010000011101000100000001110100010000000111010001000000011101000100000001110100010000000") port map( O =>C_60_S_4_out, I0 =>  C_60_S_4_L_0_out, I1 =>  C_60_S_4_L_1_out, I2 =>  C_60_S_4_L_2_out, I3 =>  C_60_S_4_L_3_out, I4 =>  C_60_S_4_L_4_out, I5 =>  C_60_S_4_L_5_out, I6 =>  C_60_S_4_L_6_out, I7 =>  C_60_S_4_L_7_out); 

C_60_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_60_out, I0 =>  C_60_S_0_out, I1 =>  C_60_S_1_out, I2 =>  C_60_S_2_out, I3 =>  C_60_S_3_out, I4 =>  C_60_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_61_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_61_S_0_out, I0 =>  C_61_S_0_L_0_out, I1 =>  C_61_S_0_L_1_out, I2 =>  C_61_S_0_L_2_out, I3 =>  C_61_S_0_L_3_out, I4 =>  C_61_S_0_L_4_out, I5 =>  C_61_S_0_L_5_out, I6 =>  C_61_S_0_L_6_out, I7 =>  C_61_S_0_L_7_out); 
C_61_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_61_S_1_out, I0 =>  C_61_S_1_L_0_out, I1 =>  C_61_S_1_L_1_out, I2 =>  C_61_S_1_L_2_out, I3 =>  C_61_S_1_L_3_out, I4 =>  C_61_S_1_L_4_out, I5 =>  C_61_S_1_L_5_out, I6 =>  C_61_S_1_L_6_out, I7 =>  C_61_S_1_L_7_out); 
C_61_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_61_S_2_out, I0 =>  C_61_S_2_L_0_out, I1 =>  C_61_S_2_L_1_out, I2 =>  C_61_S_2_L_2_out, I3 =>  C_61_S_2_L_3_out, I4 =>  C_61_S_2_L_4_out, I5 =>  C_61_S_2_L_5_out, I6 =>  C_61_S_2_L_6_out, I7 =>  C_61_S_2_L_7_out); 
C_61_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_61_S_3_out, I0 =>  C_61_S_3_L_0_out, I1 =>  C_61_S_3_L_1_out, I2 =>  C_61_S_3_L_2_out, I3 =>  C_61_S_3_L_3_out, I4 =>  C_61_S_3_L_4_out, I5 =>  C_61_S_3_L_5_out, I6 =>  C_61_S_3_L_6_out, I7 =>  C_61_S_3_L_7_out); 
C_61_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_61_S_4_out, I0 =>  C_61_S_4_L_0_out, I1 =>  C_61_S_4_L_1_out, I2 =>  C_61_S_4_L_2_out, I3 =>  C_61_S_4_L_3_out, I4 =>  C_61_S_4_L_4_out, I5 =>  C_61_S_4_L_5_out, I6 =>  C_61_S_4_L_6_out, I7 =>  C_61_S_4_L_7_out); 

C_61_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_61_out, I0 =>  C_61_S_0_out, I1 =>  C_61_S_1_out, I2 =>  C_61_S_2_out, I3 =>  C_61_S_3_out, I4 =>  C_61_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_62_S_0_inst : LUT8 generic map(INIT => "1111111011101010111011101110101011101110111010101110101010101000111010101010100011101010101010001110101010101000101010001010100011101010111010101110101010101000111010101010100011101010101010001110101010101000101010001000100010101000100010001010100010000000") port map( O =>C_62_S_0_out, I0 =>  C_62_S_0_L_0_out, I1 =>  C_62_S_0_L_1_out, I2 =>  C_62_S_0_L_2_out, I3 =>  C_62_S_0_L_3_out, I4 =>  C_62_S_0_L_4_out, I5 =>  C_62_S_0_L_5_out, I6 =>  C_62_S_0_L_6_out, I7 =>  C_62_S_0_L_7_out); 
C_62_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010100011101010101010101010101010101010101010101010101010101010101010001010101010101010101010101010100010101010101010001010100010000000") port map( O =>C_62_S_1_out, I0 =>  C_62_S_1_L_0_out, I1 =>  C_62_S_1_L_1_out, I2 =>  C_62_S_1_L_2_out, I3 =>  C_62_S_1_L_3_out, I4 =>  C_62_S_1_L_4_out, I5 =>  C_62_S_1_L_5_out, I6 =>  C_62_S_1_L_6_out, I7 =>  C_62_S_1_L_7_out); 
C_62_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111111110110011111111111011001110111011001000111111101110100011101000100000001110100010000000100010000000000011111111111011101111111011101000111111101110100011101000100000001110110010001000110010000000000011001000000000001000000000000000") port map( O =>C_62_S_2_out, I0 =>  C_62_S_2_L_0_out, I1 =>  C_62_S_2_L_1_out, I2 =>  C_62_S_2_L_2_out, I3 =>  C_62_S_2_L_3_out, I4 =>  C_62_S_2_L_4_out, I5 =>  C_62_S_2_L_5_out, I6 =>  C_62_S_2_L_6_out, I7 =>  C_62_S_2_L_7_out); 
C_62_S_3_inst : LUT8 generic map(INIT => "1111111011101110111111101110100011111110111010001110100010000000111111101110100011101100110010001110100010001000111010001000000011111110111010001110111011101000111011001100100011101000100000001111111011101000111010001000000011101000100000001000100010000000") port map( O =>C_62_S_3_out, I0 =>  C_62_S_3_L_0_out, I1 =>  C_62_S_3_L_1_out, I2 =>  C_62_S_3_L_2_out, I3 =>  C_62_S_3_L_3_out, I4 =>  C_62_S_3_L_4_out, I5 =>  C_62_S_3_L_5_out, I6 =>  C_62_S_3_L_6_out, I7 =>  C_62_S_3_L_7_out); 
C_62_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111011101110100010001000111111101110111011101010111010001110101011101000100010001000000011111110111011101110100010101000111010001010100010001000100000001110111011101000100010001000000010001000100000001000000000000000") port map( O =>C_62_S_4_out, I0 =>  C_62_S_4_L_0_out, I1 =>  C_62_S_4_L_1_out, I2 =>  C_62_S_4_L_2_out, I3 =>  C_62_S_4_L_3_out, I4 =>  C_62_S_4_L_4_out, I5 =>  C_62_S_4_L_5_out, I6 =>  C_62_S_4_L_6_out, I7 =>  C_62_S_4_L_7_out); 

C_62_inst : LUT8 generic map(INIT => "1110101011101000111010001010100011101010111010001110100010101000111010101110100011101000101010001110101011101000111010001010100011101010111010001110100010101000111010101110100011101000101010001110101011101000111010001010100011101010111010001110100010101000") port map( O =>C_62_out, I0 =>  C_62_S_0_out, I1 =>  C_62_S_1_out, I2 =>  C_62_S_2_out, I3 =>  C_62_S_3_out, I4 =>  C_62_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_63_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111111111111101111111011101000111111101110100011101000100000001110100010000000100000000000000011111111111111101111111011101000111111101110100011101000100000001110100010000000100000000000000011101000100000001000000000000000") port map( O =>C_63_S_0_out, I0 =>  C_63_S_0_L_0_out, I1 =>  C_63_S_0_L_1_out, I2 =>  C_63_S_0_L_2_out, I3 =>  C_63_S_0_L_3_out, I4 =>  C_63_S_0_L_4_out, I5 =>  C_63_S_0_L_5_out, I6 =>  C_63_S_0_L_6_out, I7 =>  C_63_S_0_L_7_out); 
C_63_S_1_inst : LUT8 generic map(INIT => "1111111111111010111111101110100011111110111010001111111010100000111111101110100011111110101010001111101010000000111010001000000011111110111010001111111010100000111010101000000011101000100000001111101010000000111010001000000011101000100000001010000000000000") port map( O =>C_63_S_1_out, I0 =>  C_63_S_1_L_0_out, I1 =>  C_63_S_1_L_1_out, I2 =>  C_63_S_1_L_2_out, I3 =>  C_63_S_1_L_3_out, I4 =>  C_63_S_1_L_4_out, I5 =>  C_63_S_1_L_5_out, I6 =>  C_63_S_1_L_6_out, I7 =>  C_63_S_1_L_7_out); 
C_63_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001111101010100000111111101110100011111010101000001111101010100000111010001000000011111110111010001111101010100000111110101010000011101000100000001111101010100000111010001000000011101000100000001000000000000000") port map( O =>C_63_S_2_out, I0 =>  C_63_S_2_L_0_out, I1 =>  C_63_S_2_L_1_out, I2 =>  C_63_S_2_L_2_out, I3 =>  C_63_S_2_L_3_out, I4 =>  C_63_S_2_L_4_out, I5 =>  C_63_S_2_L_5_out, I6 =>  C_63_S_2_L_6_out, I7 =>  C_63_S_2_L_7_out); 
C_63_S_3_inst : LUT8 generic map(INIT => "1111111111111010111111101110100011111110111010001111101010100000111111101110100011111110101000001111111011101000111010001000000011111110111010001110100010000000111110101000000011101000100000001111101010100000111010001000000011101000100000001010000000000000") port map( O =>C_63_S_3_out, I0 =>  C_63_S_3_L_0_out, I1 =>  C_63_S_3_L_1_out, I2 =>  C_63_S_3_L_2_out, I3 =>  C_63_S_3_L_3_out, I4 =>  C_63_S_3_L_4_out, I5 =>  C_63_S_3_L_5_out, I6 =>  C_63_S_3_L_6_out, I7 =>  C_63_S_3_L_7_out); 
C_63_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011101000100000001111111011101000100000000000000011111111111111101110100010000000111111101110100010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_63_S_4_out, I0 =>  C_63_S_4_L_0_out, I1 =>  C_63_S_4_L_1_out, I2 =>  C_63_S_4_L_2_out, I3 =>  C_63_S_4_L_3_out, I4 =>  C_63_S_4_L_4_out, I5 =>  C_63_S_4_L_5_out, I6 =>  C_63_S_4_L_6_out, I7 =>  C_63_S_4_L_7_out); 

C_63_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_63_out, I0 =>  C_63_S_0_out, I1 =>  C_63_S_1_out, I2 =>  C_63_S_2_out, I3 =>  C_63_S_3_out, I4 =>  C_63_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_64_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_64_S_0_out, I0 =>  C_64_S_0_L_0_out, I1 =>  C_64_S_0_L_1_out, I2 =>  C_64_S_0_L_2_out, I3 =>  C_64_S_0_L_3_out, I4 =>  C_64_S_0_L_4_out, I5 =>  C_64_S_0_L_5_out, I6 =>  C_64_S_0_L_6_out, I7 =>  C_64_S_0_L_7_out); 
C_64_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_64_S_1_out, I0 =>  C_64_S_1_L_0_out, I1 =>  C_64_S_1_L_1_out, I2 =>  C_64_S_1_L_2_out, I3 =>  C_64_S_1_L_3_out, I4 =>  C_64_S_1_L_4_out, I5 =>  C_64_S_1_L_5_out, I6 =>  C_64_S_1_L_6_out, I7 =>  C_64_S_1_L_7_out); 
C_64_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_64_S_2_out, I0 =>  C_64_S_2_L_0_out, I1 =>  C_64_S_2_L_1_out, I2 =>  C_64_S_2_L_2_out, I3 =>  C_64_S_2_L_3_out, I4 =>  C_64_S_2_L_4_out, I5 =>  C_64_S_2_L_5_out, I6 =>  C_64_S_2_L_6_out, I7 =>  C_64_S_2_L_7_out); 
C_64_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_64_S_3_out, I0 =>  C_64_S_3_L_0_out, I1 =>  C_64_S_3_L_1_out, I2 =>  C_64_S_3_L_2_out, I3 =>  C_64_S_3_L_3_out, I4 =>  C_64_S_3_L_4_out, I5 =>  C_64_S_3_L_5_out, I6 =>  C_64_S_3_L_6_out, I7 =>  C_64_S_3_L_7_out); 
C_64_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_64_S_4_out, I0 =>  C_64_S_4_L_0_out, I1 =>  C_64_S_4_L_1_out, I2 =>  C_64_S_4_L_2_out, I3 =>  C_64_S_4_L_3_out, I4 =>  C_64_S_4_L_4_out, I5 =>  C_64_S_4_L_5_out, I6 =>  C_64_S_4_L_6_out, I7 =>  C_64_S_4_L_7_out); 

C_64_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_64_out, I0 =>  C_64_S_0_out, I1 =>  C_64_S_1_out, I2 =>  C_64_S_2_out, I3 =>  C_64_S_3_out, I4 =>  C_64_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_65_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111001111110011000000111111111111110011111100110000001110100011000000100000000000000011111111111111101111110011101000111111001100000011000000000000001111110011000000110000000000000010000000000000000000000000000000") port map( O =>C_65_S_0_out, I0 =>  C_65_S_0_L_0_out, I1 =>  C_65_S_0_L_1_out, I2 =>  C_65_S_0_L_2_out, I3 =>  C_65_S_0_L_3_out, I4 =>  C_65_S_0_L_4_out, I5 =>  C_65_S_0_L_5_out, I6 =>  C_65_S_0_L_6_out, I7 =>  C_65_S_0_L_7_out); 
C_65_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111110111010001111111011001000111010000000000011111111111010001110110010000000111010001000000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_65_S_1_out, I0 =>  C_65_S_1_L_0_out, I1 =>  C_65_S_1_L_1_out, I2 =>  C_65_S_1_L_2_out, I3 =>  C_65_S_1_L_3_out, I4 =>  C_65_S_1_L_4_out, I5 =>  C_65_S_1_L_5_out, I6 =>  C_65_S_1_L_6_out, I7 =>  C_65_S_1_L_7_out); 
C_65_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111111111011111110111010001111111010100000111010000000000011111111111010001111101010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_65_S_2_out, I0 =>  C_65_S_2_L_0_out, I1 =>  C_65_S_2_L_1_out, I2 =>  C_65_S_2_L_2_out, I3 =>  C_65_S_2_L_3_out, I4 =>  C_65_S_2_L_4_out, I5 =>  C_65_S_2_L_5_out, I6 =>  C_65_S_2_L_6_out, I7 =>  C_65_S_2_L_7_out); 
C_65_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111010001111111011101000111111111110100011111110111010001110100010000000101000000000000011111111111110101111111011101000111010001000000011101000000000001110100010000000111010000000000010000000000000000000000000000000") port map( O =>C_65_S_3_out, I0 =>  C_65_S_3_L_0_out, I1 =>  C_65_S_3_L_1_out, I2 =>  C_65_S_3_L_2_out, I3 =>  C_65_S_3_L_3_out, I4 =>  C_65_S_3_L_4_out, I5 =>  C_65_S_3_L_5_out, I6 =>  C_65_S_3_L_6_out, I7 =>  C_65_S_3_L_7_out); 
C_65_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011100000111111111111111011111110111010001111111010000000100000000000000011111111111111101111111010000000111010001000000010000000000000001111100010000000100000000000000010000000000000000000000000000000") port map( O =>C_65_S_4_out, I0 =>  C_65_S_4_L_0_out, I1 =>  C_65_S_4_L_1_out, I2 =>  C_65_S_4_L_2_out, I3 =>  C_65_S_4_L_3_out, I4 =>  C_65_S_4_L_4_out, I5 =>  C_65_S_4_L_5_out, I6 =>  C_65_S_4_L_6_out, I7 =>  C_65_S_4_L_7_out); 

C_65_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_65_out, I0 =>  C_65_S_0_out, I1 =>  C_65_S_1_out, I2 =>  C_65_S_2_out, I3 =>  C_65_S_3_out, I4 =>  C_65_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_66_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_66_S_0_out, I0 =>  C_66_S_0_L_0_out, I1 =>  C_66_S_0_L_1_out, I2 =>  C_66_S_0_L_2_out, I3 =>  C_66_S_0_L_3_out, I4 =>  C_66_S_0_L_4_out, I5 =>  C_66_S_0_L_5_out, I6 =>  C_66_S_0_L_6_out, I7 =>  C_66_S_0_L_7_out); 
C_66_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_66_S_1_out, I0 =>  C_66_S_1_L_0_out, I1 =>  C_66_S_1_L_1_out, I2 =>  C_66_S_1_L_2_out, I3 =>  C_66_S_1_L_3_out, I4 =>  C_66_S_1_L_4_out, I5 =>  C_66_S_1_L_5_out, I6 =>  C_66_S_1_L_6_out, I7 =>  C_66_S_1_L_7_out); 
C_66_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_66_S_2_out, I0 =>  C_66_S_2_L_0_out, I1 =>  C_66_S_2_L_1_out, I2 =>  C_66_S_2_L_2_out, I3 =>  C_66_S_2_L_3_out, I4 =>  C_66_S_2_L_4_out, I5 =>  C_66_S_2_L_5_out, I6 =>  C_66_S_2_L_6_out, I7 =>  C_66_S_2_L_7_out); 
C_66_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_66_S_3_out, I0 =>  C_66_S_3_L_0_out, I1 =>  C_66_S_3_L_1_out, I2 =>  C_66_S_3_L_2_out, I3 =>  C_66_S_3_L_3_out, I4 =>  C_66_S_3_L_4_out, I5 =>  C_66_S_3_L_5_out, I6 =>  C_66_S_3_L_6_out, I7 =>  C_66_S_3_L_7_out); 
C_66_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_66_S_4_out, I0 =>  C_66_S_4_L_0_out, I1 =>  C_66_S_4_L_1_out, I2 =>  C_66_S_4_L_2_out, I3 =>  C_66_S_4_L_3_out, I4 =>  C_66_S_4_L_4_out, I5 =>  C_66_S_4_L_5_out, I6 =>  C_66_S_4_L_6_out, I7 =>  C_66_S_4_L_7_out); 

C_66_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_66_out, I0 =>  C_66_S_0_out, I1 =>  C_66_S_1_out, I2 =>  C_66_S_2_out, I3 =>  C_66_S_3_out, I4 =>  C_66_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_67_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011100000111111111111111011111110101000001111100010000000100000000000000011111111111111101111111011100000111110101000000010000000000000001111100010000000100000000000000010000000000000000000000000000000") port map( O =>C_67_S_0_out, I0 =>  C_67_S_0_L_0_out, I1 =>  C_67_S_0_L_1_out, I2 =>  C_67_S_0_L_2_out, I3 =>  C_67_S_0_L_3_out, I4 =>  C_67_S_0_L_4_out, I5 =>  C_67_S_0_L_5_out, I6 =>  C_67_S_0_L_6_out, I7 =>  C_67_S_0_L_7_out); 
C_67_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111010000000111111111111111011111110111000001111111010000000101000000000000011111111111110101111111010000000111110001000000010000000000000001111111010000000100000000000000010000000000000000000000000000000") port map( O =>C_67_S_1_out, I0 =>  C_67_S_1_L_0_out, I1 =>  C_67_S_1_L_1_out, I2 =>  C_67_S_1_L_2_out, I3 =>  C_67_S_1_L_3_out, I4 =>  C_67_S_1_L_4_out, I5 =>  C_67_S_1_L_5_out, I6 =>  C_67_S_1_L_6_out, I7 =>  C_67_S_1_L_7_out); 
C_67_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111110101111111010000000111111111111111011111110111000001111100010000000100000000000000011111111111111101111111011100000111110001000000010000000000000001111111010000000101000000000000010000000000000000000000000000000") port map( O =>C_67_S_2_out, I0 =>  C_67_S_2_L_0_out, I1 =>  C_67_S_2_L_1_out, I2 =>  C_67_S_2_L_2_out, I3 =>  C_67_S_2_L_3_out, I4 =>  C_67_S_2_L_4_out, I5 =>  C_67_S_2_L_5_out, I6 =>  C_67_S_2_L_6_out, I7 =>  C_67_S_2_L_7_out); 
C_67_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111110001111100010000000111111111111111011111110111000001111100010000000100000000000000011111111111111101111111011100000111110001000000010000000000000001111111011100000111000000000000010000000000000000000000000000000") port map( O =>C_67_S_3_out, I0 =>  C_67_S_3_L_0_out, I1 =>  C_67_S_3_L_1_out, I2 =>  C_67_S_3_L_2_out, I3 =>  C_67_S_3_L_3_out, I4 =>  C_67_S_3_L_4_out, I5 =>  C_67_S_3_L_5_out, I6 =>  C_67_S_3_L_6_out, I7 =>  C_67_S_3_L_7_out); 
C_67_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111110011101000111111111111111011111100111010001111110011101000110000001000000011111110111111001110100011000000111010001100000010000000000000001110100011000000100000000000000010000000000000000000000000000000") port map( O =>C_67_S_4_out, I0 =>  C_67_S_4_L_0_out, I1 =>  C_67_S_4_L_1_out, I2 =>  C_67_S_4_L_2_out, I3 =>  C_67_S_4_L_3_out, I4 =>  C_67_S_4_L_4_out, I5 =>  C_67_S_4_L_5_out, I6 =>  C_67_S_4_L_6_out, I7 =>  C_67_S_4_L_7_out); 

C_67_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_67_out, I0 =>  C_67_S_0_out, I1 =>  C_67_S_1_out, I2 =>  C_67_S_2_out, I3 =>  C_67_S_3_out, I4 =>  C_67_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_68_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111001111110011000000111111111111110011111100110000001110100011000000100000000000000011111111111111101111110011101000111111001100000011000000000000001111110011000000110000000000000010000000000000000000000000000000") port map( O =>C_68_S_0_out, I0 =>  C_68_S_0_L_0_out, I1 =>  C_68_S_0_L_1_out, I2 =>  C_68_S_0_L_2_out, I3 =>  C_68_S_0_L_3_out, I4 =>  C_68_S_0_L_4_out, I5 =>  C_68_S_0_L_5_out, I6 =>  C_68_S_0_L_6_out, I7 =>  C_68_S_0_L_7_out); 
C_68_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101110100010000000111111111111111011111110110010001111111011001000100000000000000011111111111111101110110010000000111011001000000010000000000000001111111011101000100000000000000010000000000000000000000000000000") port map( O =>C_68_S_1_out, I0 =>  C_68_S_1_L_0_out, I1 =>  C_68_S_1_L_1_out, I2 =>  C_68_S_1_L_2_out, I3 =>  C_68_S_1_L_3_out, I4 =>  C_68_S_1_L_4_out, I5 =>  C_68_S_1_L_5_out, I6 =>  C_68_S_1_L_6_out, I7 =>  C_68_S_1_L_7_out); 
C_68_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111111111100011111110101000001111100010000000101000000000000011111111111110101111111011100000111110101000000011100000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_68_S_2_out, I0 =>  C_68_S_2_L_0_out, I1 =>  C_68_S_2_L_1_out, I2 =>  C_68_S_2_L_2_out, I3 =>  C_68_S_2_L_3_out, I4 =>  C_68_S_2_L_4_out, I5 =>  C_68_S_2_L_5_out, I6 =>  C_68_S_2_L_6_out, I7 =>  C_68_S_2_L_7_out); 
C_68_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111110111010001111111011100000111111111111111011111110111010001111111010100000111010001000000011111110111010001111101010000000111010001000000010000000000000001111100010000000111010001000000010000000000000000000000000000000") port map( O =>C_68_S_3_out, I0 =>  C_68_S_3_L_0_out, I1 =>  C_68_S_3_L_1_out, I2 =>  C_68_S_3_L_2_out, I3 =>  C_68_S_3_L_3_out, I4 =>  C_68_S_3_L_4_out, I5 =>  C_68_S_3_L_5_out, I6 =>  C_68_S_3_L_6_out, I7 =>  C_68_S_3_L_7_out); 
C_68_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011100000111111111111111011111110111010001111111010000000100000000000000011111111111111101111111010000000111010001000000010000000000000001111100010000000100000000000000010000000000000000000000000000000") port map( O =>C_68_S_4_out, I0 =>  C_68_S_4_L_0_out, I1 =>  C_68_S_4_L_1_out, I2 =>  C_68_S_4_L_2_out, I3 =>  C_68_S_4_L_3_out, I4 =>  C_68_S_4_L_4_out, I5 =>  C_68_S_4_L_5_out, I6 =>  C_68_S_4_L_6_out, I7 =>  C_68_S_4_L_7_out); 

C_68_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_68_out, I0 =>  C_68_S_0_out, I1 =>  C_68_S_1_out, I2 =>  C_68_S_2_out, I3 =>  C_68_S_3_out, I4 =>  C_68_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_69_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_69_S_0_out, I0 =>  C_69_S_0_L_0_out, I1 =>  C_69_S_0_L_1_out, I2 =>  C_69_S_0_L_2_out, I3 =>  C_69_S_0_L_3_out, I4 =>  C_69_S_0_L_4_out, I5 =>  C_69_S_0_L_5_out, I6 =>  C_69_S_0_L_6_out, I7 =>  C_69_S_0_L_7_out); 
C_69_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_69_S_1_out, I0 =>  C_69_S_1_L_0_out, I1 =>  C_69_S_1_L_1_out, I2 =>  C_69_S_1_L_2_out, I3 =>  C_69_S_1_L_3_out, I4 =>  C_69_S_1_L_4_out, I5 =>  C_69_S_1_L_5_out, I6 =>  C_69_S_1_L_6_out, I7 =>  C_69_S_1_L_7_out); 
C_69_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_69_S_2_out, I0 =>  C_69_S_2_L_0_out, I1 =>  C_69_S_2_L_1_out, I2 =>  C_69_S_2_L_2_out, I3 =>  C_69_S_2_L_3_out, I4 =>  C_69_S_2_L_4_out, I5 =>  C_69_S_2_L_5_out, I6 =>  C_69_S_2_L_6_out, I7 =>  C_69_S_2_L_7_out); 
C_69_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111111111111011111110111000001111111010000000100000000000000011111111111111101111111010000000111110001000000010000000000000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_69_S_3_out, I0 =>  C_69_S_3_L_0_out, I1 =>  C_69_S_3_L_1_out, I2 =>  C_69_S_3_L_2_out, I3 =>  C_69_S_3_L_3_out, I4 =>  C_69_S_3_L_4_out, I5 =>  C_69_S_3_L_5_out, I6 =>  C_69_S_3_L_6_out, I7 =>  C_69_S_3_L_7_out); 
C_69_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_69_S_4_out, I0 =>  C_69_S_4_L_0_out, I1 =>  C_69_S_4_L_1_out, I2 =>  C_69_S_4_L_2_out, I3 =>  C_69_S_4_L_3_out, I4 =>  C_69_S_4_L_4_out, I5 =>  C_69_S_4_L_5_out, I6 =>  C_69_S_4_L_6_out, I7 =>  C_69_S_4_L_7_out); 

C_69_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_69_out, I0 =>  C_69_S_0_out, I1 =>  C_69_S_1_out, I2 =>  C_69_S_2_out, I3 =>  C_69_S_3_out, I4 =>  C_69_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_70_S_0_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_70_S_0_out, I0 =>  C_70_S_0_L_0_out, I1 =>  C_70_S_0_L_1_out, I2 =>  C_70_S_0_L_2_out, I3 =>  C_70_S_0_L_3_out, I4 =>  C_70_S_0_L_4_out, I5 =>  C_70_S_0_L_5_out, I6 =>  C_70_S_0_L_6_out, I7 =>  C_70_S_0_L_7_out); 
C_70_S_1_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_70_S_1_out, I0 =>  C_70_S_1_L_0_out, I1 =>  C_70_S_1_L_1_out, I2 =>  C_70_S_1_L_2_out, I3 =>  C_70_S_1_L_3_out, I4 =>  C_70_S_1_L_4_out, I5 =>  C_70_S_1_L_5_out, I6 =>  C_70_S_1_L_6_out, I7 =>  C_70_S_1_L_7_out); 
C_70_S_2_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_70_S_2_out, I0 =>  C_70_S_2_L_0_out, I1 =>  C_70_S_2_L_1_out, I2 =>  C_70_S_2_L_2_out, I3 =>  C_70_S_2_L_3_out, I4 =>  C_70_S_2_L_4_out, I5 =>  C_70_S_2_L_5_out, I6 =>  C_70_S_2_L_6_out, I7 =>  C_70_S_2_L_7_out); 
C_70_S_3_inst : LUT8 generic map(INIT => "1111111111101110111111101110100011111110111010001110111010001000111011101110100011101110100010001110111010001000111010001000000011111110111010001110111010001000111011101000100011101000100010001110111010001000111010001000000011101000100000001000100000000000") port map( O =>C_70_S_3_out, I0 =>  C_70_S_3_L_0_out, I1 =>  C_70_S_3_L_1_out, I2 =>  C_70_S_3_L_2_out, I3 =>  C_70_S_3_L_3_out, I4 =>  C_70_S_3_L_4_out, I5 =>  C_70_S_3_L_5_out, I6 =>  C_70_S_3_L_6_out, I7 =>  C_70_S_3_L_7_out); 
C_70_S_4_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_70_S_4_out, I0 =>  C_70_S_4_L_0_out, I1 =>  C_70_S_4_L_1_out, I2 =>  C_70_S_4_L_2_out, I3 =>  C_70_S_4_L_3_out, I4 =>  C_70_S_4_L_4_out, I5 =>  C_70_S_4_L_5_out, I6 =>  C_70_S_4_L_6_out, I7 =>  C_70_S_4_L_7_out); 

C_70_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_70_out, I0 =>  C_70_S_0_out, I1 =>  C_70_S_1_out, I2 =>  C_70_S_2_out, I3 =>  C_70_S_3_out, I4 =>  C_70_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_71_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001111101010000000111111101110100011111110100000001111111010000000111010001000000011111110111010001111111010000000111111101000000011101000100000001111111010100000111010001000000011101000100000001000000000000000") port map( O =>C_71_S_0_out, I0 =>  C_71_S_0_L_0_out, I1 =>  C_71_S_0_L_1_out, I2 =>  C_71_S_0_L_2_out, I3 =>  C_71_S_0_L_3_out, I4 =>  C_71_S_0_L_4_out, I5 =>  C_71_S_0_L_5_out, I6 =>  C_71_S_0_L_6_out, I7 =>  C_71_S_0_L_7_out); 
C_71_S_1_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_71_S_1_out, I0 =>  C_71_S_1_L_0_out, I1 =>  C_71_S_1_L_1_out, I2 =>  C_71_S_1_L_2_out, I3 =>  C_71_S_1_L_3_out, I4 =>  C_71_S_1_L_4_out, I5 =>  C_71_S_1_L_5_out, I6 =>  C_71_S_1_L_6_out, I7 =>  C_71_S_1_L_7_out); 
C_71_S_2_inst : LUT8 generic map(INIT => "1111111111111000111111101110100011111110111010001111111010100000111111101110100011111000100000001111101010000000111010001000000011111110111010001111111010100000111111101110000011101000100000001111101010000000111010001000000011101000100000001110000000000000") port map( O =>C_71_S_2_out, I0 =>  C_71_S_2_L_0_out, I1 =>  C_71_S_2_L_1_out, I2 =>  C_71_S_2_L_2_out, I3 =>  C_71_S_2_L_3_out, I4 =>  C_71_S_2_L_4_out, I5 =>  C_71_S_2_L_5_out, I6 =>  C_71_S_2_L_6_out, I7 =>  C_71_S_2_L_7_out); 
C_71_S_3_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_71_S_3_out, I0 =>  C_71_S_3_L_0_out, I1 =>  C_71_S_3_L_1_out, I2 =>  C_71_S_3_L_2_out, I3 =>  C_71_S_3_L_3_out, I4 =>  C_71_S_3_L_4_out, I5 =>  C_71_S_3_L_5_out, I6 =>  C_71_S_3_L_6_out, I7 =>  C_71_S_3_L_7_out); 
C_71_S_4_inst : LUT8 generic map(INIT => "1111111111101110111111101110100011111110111010001111111010001000111111101110100011111110100010001110111010000000111010001000000011111110111010001111111010001000111011101000000011101000100000001110111010000000111010001000000011101000100000001000100000000000") port map( O =>C_71_S_4_out, I0 =>  C_71_S_4_L_0_out, I1 =>  C_71_S_4_L_1_out, I2 =>  C_71_S_4_L_2_out, I3 =>  C_71_S_4_L_3_out, I4 =>  C_71_S_4_L_4_out, I5 =>  C_71_S_4_L_5_out, I6 =>  C_71_S_4_L_6_out, I7 =>  C_71_S_4_L_7_out); 

C_71_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_71_out, I0 =>  C_71_S_0_out, I1 =>  C_71_S_1_out, I2 =>  C_71_S_2_out, I3 =>  C_71_S_3_out, I4 =>  C_71_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_72_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101110100011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100011101000101010001010100010000000") port map( O =>C_72_S_0_out, I0 =>  C_72_S_0_L_0_out, I1 =>  C_72_S_0_L_1_out, I2 =>  C_72_S_0_L_2_out, I3 =>  C_72_S_0_L_3_out, I4 =>  C_72_S_0_L_4_out, I5 =>  C_72_S_0_L_5_out, I6 =>  C_72_S_0_L_6_out, I7 =>  C_72_S_0_L_7_out); 
C_72_S_1_inst : LUT8 generic map(INIT => "1111111011101010111010101110100011101110111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001000100011101000101010001010100010000000") port map( O =>C_72_S_1_out, I0 =>  C_72_S_1_L_0_out, I1 =>  C_72_S_1_L_1_out, I2 =>  C_72_S_1_L_2_out, I3 =>  C_72_S_1_L_3_out, I4 =>  C_72_S_1_L_4_out, I5 =>  C_72_S_1_L_5_out, I6 =>  C_72_S_1_L_6_out, I7 =>  C_72_S_1_L_7_out); 
C_72_S_2_inst : LUT8 generic map(INIT => "1111111011101010111011101110101011101010111010101110101010101000111010101110101011101010101010001110101010101000101010001010100011101010111010101110101010101000111010101010100010101000101010001110101010101000101010001010100010101000100010001010100010000000") port map( O =>C_72_S_2_out, I0 =>  C_72_S_2_L_0_out, I1 =>  C_72_S_2_L_1_out, I2 =>  C_72_S_2_L_2_out, I3 =>  C_72_S_2_L_3_out, I4 =>  C_72_S_2_L_4_out, I5 =>  C_72_S_2_L_5_out, I6 =>  C_72_S_2_L_6_out, I7 =>  C_72_S_2_L_7_out); 
C_72_S_3_inst : LUT8 generic map(INIT => "1111111011101110111111101110100011111110111010001110111011101000111111101110100011101010101010001110111011101000111010001000000011111110111010001110100010001000111010101010100011101000100000001110100010001000111010001000000011101000100000001000100010000000") port map( O =>C_72_S_3_out, I0 =>  C_72_S_3_L_0_out, I1 =>  C_72_S_3_L_1_out, I2 =>  C_72_S_3_L_2_out, I3 =>  C_72_S_3_L_3_out, I4 =>  C_72_S_3_L_4_out, I5 =>  C_72_S_3_L_5_out, I6 =>  C_72_S_3_L_6_out, I7 =>  C_72_S_3_L_7_out); 
C_72_S_4_inst : LUT8 generic map(INIT => "1111111011101110111011101110100011101110111010001110100011101000111011101110100011101000111010001110100011101000111010001000100011101110111010001110100011101000111010001110100011101000100010001110100011101000111010001000100011101000100010001000100010000000") port map( O =>C_72_S_4_out, I0 =>  C_72_S_4_L_0_out, I1 =>  C_72_S_4_L_1_out, I2 =>  C_72_S_4_L_2_out, I3 =>  C_72_S_4_L_3_out, I4 =>  C_72_S_4_L_4_out, I5 =>  C_72_S_4_L_5_out, I6 =>  C_72_S_4_L_6_out, I7 =>  C_72_S_4_L_7_out); 

C_72_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_72_out, I0 =>  C_72_S_0_out, I1 =>  C_72_S_1_out, I2 =>  C_72_S_2_out, I3 =>  C_72_S_3_out, I4 =>  C_72_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_73_S_0_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001000000010000000") port map( O =>C_73_S_0_out, I0 =>  C_73_S_0_L_0_out, I1 =>  C_73_S_0_L_1_out, I2 =>  C_73_S_0_L_2_out, I3 =>  C_73_S_0_L_3_out, I4 =>  C_73_S_0_L_4_out, I5 =>  C_73_S_0_L_5_out, I6 =>  C_73_S_0_L_6_out, I7 =>  C_73_S_0_L_7_out); 
C_73_S_1_inst : LUT8 generic map(INIT => "1111111011111110111011101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100010001000000010000000") port map( O =>C_73_S_1_out, I0 =>  C_73_S_1_L_0_out, I1 =>  C_73_S_1_L_1_out, I2 =>  C_73_S_1_L_2_out, I3 =>  C_73_S_1_L_3_out, I4 =>  C_73_S_1_L_4_out, I5 =>  C_73_S_1_L_5_out, I6 =>  C_73_S_1_L_6_out, I7 =>  C_73_S_1_L_7_out); 
C_73_S_2_inst : LUT8 generic map(INIT => "1111111011101110111111101110100011101110111010001110100010101000111011101110100011101000101010001110100010001000101010001000000011111110111010101110111011101000111010101110100011101000100010001110101011101000111010001000100011101000100000001000100010000000") port map( O =>C_73_S_2_out, I0 =>  C_73_S_2_L_0_out, I1 =>  C_73_S_2_L_1_out, I2 =>  C_73_S_2_L_2_out, I3 =>  C_73_S_2_L_3_out, I4 =>  C_73_S_2_L_4_out, I5 =>  C_73_S_2_L_5_out, I6 =>  C_73_S_2_L_6_out, I7 =>  C_73_S_2_L_7_out); 
C_73_S_3_inst : LUT8 generic map(INIT => "1111111011111010111110101110100011111010111010001110100011100000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001111100011101000111010001010000011101000101000001010000010000000") port map( O =>C_73_S_3_out, I0 =>  C_73_S_3_L_0_out, I1 =>  C_73_S_3_L_1_out, I2 =>  C_73_S_3_L_2_out, I3 =>  C_73_S_3_L_3_out, I4 =>  C_73_S_3_L_4_out, I5 =>  C_73_S_3_L_5_out, I6 =>  C_73_S_3_L_6_out, I7 =>  C_73_S_3_L_7_out); 
C_73_S_4_inst : LUT8 generic map(INIT => "1111111011111110111110101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000101000001000000010000000") port map( O =>C_73_S_4_out, I0 =>  C_73_S_4_L_0_out, I1 =>  C_73_S_4_L_1_out, I2 =>  C_73_S_4_L_2_out, I3 =>  C_73_S_4_L_3_out, I4 =>  C_73_S_4_L_4_out, I5 =>  C_73_S_4_L_5_out, I6 =>  C_73_S_4_L_6_out, I7 =>  C_73_S_4_L_7_out); 

C_73_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_73_out, I0 =>  C_73_S_0_out, I1 =>  C_73_S_1_out, I2 =>  C_73_S_2_out, I3 =>  C_73_S_3_out, I4 =>  C_73_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_74_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_74_S_0_out, I0 =>  C_74_S_0_L_0_out, I1 =>  C_74_S_0_L_1_out, I2 =>  C_74_S_0_L_2_out, I3 =>  C_74_S_0_L_3_out, I4 =>  C_74_S_0_L_4_out, I5 =>  C_74_S_0_L_5_out, I6 =>  C_74_S_0_L_6_out, I7 =>  C_74_S_0_L_7_out); 
C_74_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_74_S_1_out, I0 =>  C_74_S_1_L_0_out, I1 =>  C_74_S_1_L_1_out, I2 =>  C_74_S_1_L_2_out, I3 =>  C_74_S_1_L_3_out, I4 =>  C_74_S_1_L_4_out, I5 =>  C_74_S_1_L_5_out, I6 =>  C_74_S_1_L_6_out, I7 =>  C_74_S_1_L_7_out); 
C_74_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_74_S_2_out, I0 =>  C_74_S_2_L_0_out, I1 =>  C_74_S_2_L_1_out, I2 =>  C_74_S_2_L_2_out, I3 =>  C_74_S_2_L_3_out, I4 =>  C_74_S_2_L_4_out, I5 =>  C_74_S_2_L_5_out, I6 =>  C_74_S_2_L_6_out, I7 =>  C_74_S_2_L_7_out); 
C_74_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_74_S_3_out, I0 =>  C_74_S_3_L_0_out, I1 =>  C_74_S_3_L_1_out, I2 =>  C_74_S_3_L_2_out, I3 =>  C_74_S_3_L_3_out, I4 =>  C_74_S_3_L_4_out, I5 =>  C_74_S_3_L_5_out, I6 =>  C_74_S_3_L_6_out, I7 =>  C_74_S_3_L_7_out); 
C_74_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011101000100000001110100010000000100000000000000011111110111010001110100010000000111010001000000010000000000000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_74_S_4_out, I0 =>  C_74_S_4_L_0_out, I1 =>  C_74_S_4_L_1_out, I2 =>  C_74_S_4_L_2_out, I3 =>  C_74_S_4_L_3_out, I4 =>  C_74_S_4_L_4_out, I5 =>  C_74_S_4_L_5_out, I6 =>  C_74_S_4_L_6_out, I7 =>  C_74_S_4_L_7_out); 

C_74_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_74_out, I0 =>  C_74_S_0_out, I1 =>  C_74_S_1_out, I2 =>  C_74_S_2_out, I3 =>  C_74_S_3_out, I4 =>  C_74_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_75_S_0_inst : LUT8 generic map(INIT => "1111111011111110111111101111101011111110111010001111100011101000111110101110100011101000111010001110100011101000111010001000000011111110111010001110100011101000111010001110100011101000101000001110100011100000111010001000000010100000100000001000000010000000") port map( O =>C_75_S_0_out, I0 =>  C_75_S_0_L_0_out, I1 =>  C_75_S_0_L_1_out, I2 =>  C_75_S_0_L_2_out, I3 =>  C_75_S_0_L_3_out, I4 =>  C_75_S_0_L_4_out, I5 =>  C_75_S_0_L_5_out, I6 =>  C_75_S_0_L_6_out, I7 =>  C_75_S_0_L_7_out); 
C_75_S_1_inst : LUT8 generic map(INIT => "1111111011111010111110101110100011111110111010001110100011101000111110101110100011101000111010001110100011101000111010001010000011111010111010001110100011101000111010001110100011101000101000001110100011101000111010001000000011101000101000001010000010000000") port map( O =>C_75_S_1_out, I0 =>  C_75_S_1_L_0_out, I1 =>  C_75_S_1_L_1_out, I2 =>  C_75_S_1_L_2_out, I3 =>  C_75_S_1_L_3_out, I4 =>  C_75_S_1_L_4_out, I5 =>  C_75_S_1_L_5_out, I6 =>  C_75_S_1_L_6_out, I7 =>  C_75_S_1_L_7_out); 
C_75_S_2_inst : LUT8 generic map(INIT => "1111111011111110111111101110101011111110111010001110100011101000111111101110101011101000111010001110100011101000101010001000000011111110111010101110100011101000111010001110100010101000100000001110100011101000111010001000000010101000100000001000000010000000") port map( O =>C_75_S_2_out, I0 =>  C_75_S_2_L_0_out, I1 =>  C_75_S_2_L_1_out, I2 =>  C_75_S_2_L_2_out, I3 =>  C_75_S_2_L_3_out, I4 =>  C_75_S_2_L_4_out, I5 =>  C_75_S_2_L_5_out, I6 =>  C_75_S_2_L_6_out, I7 =>  C_75_S_2_L_7_out); 
C_75_S_3_inst : LUT8 generic map(INIT => "1111111011111110111111101110100011101010111010001110100010101000111111101110100011101000111010001110100010101000101010001000000011111110111010101110101011101000111010001110100011101000100000001110101011101000111010001010100011101000100000001000000010000000") port map( O =>C_75_S_3_out, I0 =>  C_75_S_3_L_0_out, I1 =>  C_75_S_3_L_1_out, I2 =>  C_75_S_3_L_2_out, I3 =>  C_75_S_3_L_3_out, I4 =>  C_75_S_3_L_4_out, I5 =>  C_75_S_3_L_5_out, I6 =>  C_75_S_3_L_6_out, I7 =>  C_75_S_3_L_7_out); 
C_75_S_4_inst : LUT8 generic map(INIT => "1111111011111010111111101110100011111110111010001110100011101000111111101110100011101000111010001110100011101000111010001010000011111010111010001110100011101000111010001110100011101000100000001110100011101000111010001000000011101000100000001010000010000000") port map( O =>C_75_S_4_out, I0 =>  C_75_S_4_L_0_out, I1 =>  C_75_S_4_L_1_out, I2 =>  C_75_S_4_L_2_out, I3 =>  C_75_S_4_L_3_out, I4 =>  C_75_S_4_L_4_out, I5 =>  C_75_S_4_L_5_out, I6 =>  C_75_S_4_L_6_out, I7 =>  C_75_S_4_L_7_out); 

C_75_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_75_out, I0 =>  C_75_S_0_out, I1 =>  C_75_S_1_out, I2 =>  C_75_S_2_out, I3 =>  C_75_S_3_out, I4 =>  C_75_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_76_S_0_inst : LUT8 generic map(INIT => "1111111011101110111011101110101011101010111010101110101010101000111011101110101011101010101010001110101010101000101010001000100011101110111010101110101010101000111010101010100010101000100010001110101010101000101010001010100010101000100010001000100010000000") port map( O =>C_76_S_0_out, I0 =>  C_76_S_0_L_0_out, I1 =>  C_76_S_0_L_1_out, I2 =>  C_76_S_0_L_2_out, I3 =>  C_76_S_0_L_3_out, I4 =>  C_76_S_0_L_4_out, I5 =>  C_76_S_0_L_5_out, I6 =>  C_76_S_0_L_6_out, I7 =>  C_76_S_0_L_7_out); 
C_76_S_1_inst : LUT8 generic map(INIT => "1111111011101010111111101110101011101010101010001110101010101000111111101010100011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100011101010100000001110101010101000111010101010100010101000100000001010100010000000") port map( O =>C_76_S_1_out, I0 =>  C_76_S_1_L_0_out, I1 =>  C_76_S_1_L_1_out, I2 =>  C_76_S_1_L_2_out, I3 =>  C_76_S_1_L_3_out, I4 =>  C_76_S_1_L_4_out, I5 =>  C_76_S_1_L_5_out, I6 =>  C_76_S_1_L_6_out, I7 =>  C_76_S_1_L_7_out); 
C_76_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111111111010001111101010000000111111111111101011111110111010001111111011101000111010001000000011111110111010001110100010000000111010001000000010100000000000001111111010100000111010000000000011101000100000001000000000000000") port map( O =>C_76_S_2_out, I0 =>  C_76_S_2_L_0_out, I1 =>  C_76_S_2_L_1_out, I2 =>  C_76_S_2_L_2_out, I3 =>  C_76_S_2_L_3_out, I4 =>  C_76_S_2_L_4_out, I5 =>  C_76_S_2_L_5_out, I6 =>  C_76_S_2_L_6_out, I7 =>  C_76_S_2_L_7_out); 
C_76_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110101011111110111010101110101010101000111111101110101011101010101010001110101010101000101010001000000011111110111010101110101010101000111010101010100010101000100000001110101010101000101010001000000010101000100000001000000000000000") port map( O =>C_76_S_3_out, I0 =>  C_76_S_3_L_0_out, I1 =>  C_76_S_3_L_1_out, I2 =>  C_76_S_3_L_2_out, I3 =>  C_76_S_3_L_3_out, I4 =>  C_76_S_3_L_4_out, I5 =>  C_76_S_3_L_5_out, I6 =>  C_76_S_3_L_6_out, I7 =>  C_76_S_3_L_7_out); 
C_76_S_4_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111011101110111011101000111111101110111011101110111010001111111011101000111010001000000011111110111010001110100010000000111010001000100010001000100000001110100010001000100010001000000010001000100000001000000000000000") port map( O =>C_76_S_4_out, I0 =>  C_76_S_4_L_0_out, I1 =>  C_76_S_4_L_1_out, I2 =>  C_76_S_4_L_2_out, I3 =>  C_76_S_4_L_3_out, I4 =>  C_76_S_4_L_4_out, I5 =>  C_76_S_4_L_5_out, I6 =>  C_76_S_4_L_6_out, I7 =>  C_76_S_4_L_7_out); 

C_76_inst : LUT8 generic map(INIT => "1110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000111011101110100011101000100010001110111011101000111010001000100011101110111010001110100010001000") port map( O =>C_76_out, I0 =>  C_76_S_0_out, I1 =>  C_76_S_1_out, I2 =>  C_76_S_2_out, I3 =>  C_76_S_3_out, I4 =>  C_76_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_77_S_0_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111111111111101110111010001000111111101110111011101000100000001111111011101000110010001000000011111110111011001110100010000000111111101110100010001000100000001110111010001000100000000000000011101000100000001000000000000000") port map( O =>C_77_S_0_out, I0 =>  C_77_S_0_L_0_out, I1 =>  C_77_S_0_L_1_out, I2 =>  C_77_S_0_L_2_out, I3 =>  C_77_S_0_L_3_out, I4 =>  C_77_S_0_L_4_out, I5 =>  C_77_S_0_L_5_out, I6 =>  C_77_S_0_L_6_out, I7 =>  C_77_S_0_L_7_out); 
C_77_S_1_inst : LUT8 generic map(INIT => "1111111111101010111111101110100011111110111010001111111010100000111111101110100011111010100000001111101010000000111010001000000011111110111010001111111010100000111111101010000011101000100000001111101010000000111010001000000011101000100000001010100000000000") port map( O =>C_77_S_1_out, I0 =>  C_77_S_1_L_0_out, I1 =>  C_77_S_1_L_1_out, I2 =>  C_77_S_1_L_2_out, I3 =>  C_77_S_1_L_3_out, I4 =>  C_77_S_1_L_4_out, I5 =>  C_77_S_1_L_5_out, I6 =>  C_77_S_1_L_6_out, I7 =>  C_77_S_1_L_7_out); 
C_77_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111001110100011111110111110001110100010000000111111101110100011101000100000001111111011101000111000001000000011111110111110001110100010000000111111101110100011101000100000001111111011101000111000001000000011101000110000001000000000000000") port map( O =>C_77_S_2_out, I0 =>  C_77_S_2_L_0_out, I1 =>  C_77_S_2_L_1_out, I2 =>  C_77_S_2_L_2_out, I3 =>  C_77_S_2_L_3_out, I4 =>  C_77_S_2_L_4_out, I5 =>  C_77_S_2_L_5_out, I6 =>  C_77_S_2_L_6_out, I7 =>  C_77_S_2_L_7_out); 
C_77_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001111111011101000111010001000000011101000100000001000000000000000") port map( O =>C_77_S_3_out, I0 =>  C_77_S_3_L_0_out, I1 =>  C_77_S_3_L_1_out, I2 =>  C_77_S_3_L_2_out, I3 =>  C_77_S_3_L_3_out, I4 =>  C_77_S_3_L_4_out, I5 =>  C_77_S_3_L_5_out, I6 =>  C_77_S_3_L_6_out, I7 =>  C_77_S_3_L_7_out); 
C_77_S_4_inst : LUT8 generic map(INIT => "1111111111101110111111101110100011111110111010001110100010000000111111101110100011111110111010001110100010000000111010001000000011111110111010001111111011101000111010001000000011101000100000001111111011101000111010001000000011101000100000001000100000000000") port map( O =>C_77_S_4_out, I0 =>  C_77_S_4_L_0_out, I1 =>  C_77_S_4_L_1_out, I2 =>  C_77_S_4_L_2_out, I3 =>  C_77_S_4_L_3_out, I4 =>  C_77_S_4_L_4_out, I5 =>  C_77_S_4_L_5_out, I6 =>  C_77_S_4_L_6_out, I7 =>  C_77_S_4_L_7_out); 

C_77_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_77_out, I0 =>  C_77_S_0_out, I1 =>  C_77_S_1_out, I2 =>  C_77_S_2_out, I3 =>  C_77_S_3_out, I4 =>  C_77_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_78_S_0_inst : LUT8 generic map(INIT => "1111111011101010111010101010101011101010101010101010101010101000111010101010101010101010101010001110101010101010101010001010100011101010111010101010101010101000111010101010101010101010101010001110101010101010101010101010100010101010101010001010100010000000") port map( O =>C_78_S_0_out, I0 =>  C_78_S_0_L_0_out, I1 =>  C_78_S_0_L_1_out, I2 =>  C_78_S_0_L_2_out, I3 =>  C_78_S_0_L_3_out, I4 =>  C_78_S_0_L_4_out, I5 =>  C_78_S_0_L_5_out, I6 =>  C_78_S_0_L_6_out, I7 =>  C_78_S_0_L_7_out); 
C_78_S_1_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010101000111111101110101011101010111010001110100010101000101010001000000011111110111010101110101011101000111010001010100010101000100000001110101011101000111010001000000011101000100000001000000000000000") port map( O =>C_78_S_1_out, I0 =>  C_78_S_1_L_0_out, I1 =>  C_78_S_1_L_1_out, I2 =>  C_78_S_1_L_2_out, I3 =>  C_78_S_1_L_3_out, I4 =>  C_78_S_1_L_4_out, I5 =>  C_78_S_1_L_5_out, I6 =>  C_78_S_1_L_6_out, I7 =>  C_78_S_1_L_7_out); 
C_78_S_2_inst : LUT8 generic map(INIT => "1111111111111110111111101110100011111110111010001110101010100000111111101110100011101010101000001111101010100000101010001000000011111110111010101111101010100000111110101010100011101000100000001111101010101000111010001000000011101000100000001000000000000000") port map( O =>C_78_S_2_out, I0 =>  C_78_S_2_L_0_out, I1 =>  C_78_S_2_L_1_out, I2 =>  C_78_S_2_L_2_out, I3 =>  C_78_S_2_L_3_out, I4 =>  C_78_S_2_L_4_out, I5 =>  C_78_S_2_L_5_out, I6 =>  C_78_S_2_L_6_out, I7 =>  C_78_S_2_L_7_out); 
C_78_S_3_inst : LUT8 generic map(INIT => "1111111111111110111111101110111011111110111111101110111011101000111111101110111011101010111010001110111011101000111010001000000011111110111010001110100010001000111010001010100010001000100000001110100010001000100000001000000010001000100000001000000000000000") port map( O =>C_78_S_3_out, I0 =>  C_78_S_3_L_0_out, I1 =>  C_78_S_3_L_1_out, I2 =>  C_78_S_3_L_2_out, I3 =>  C_78_S_3_L_3_out, I4 =>  C_78_S_3_L_4_out, I5 =>  C_78_S_3_L_5_out, I6 =>  C_78_S_3_L_6_out, I7 =>  C_78_S_3_L_7_out); 
C_78_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111110101111111010101000111111111110101011111010101010001110101010100000101010000000000011111111111010101111101010101000111010101010000010101000000000001110101010000000101000000000000010000000000000000000000000000000") port map( O =>C_78_S_4_out, I0 =>  C_78_S_4_L_0_out, I1 =>  C_78_S_4_L_1_out, I2 =>  C_78_S_4_L_2_out, I3 =>  C_78_S_4_L_3_out, I4 =>  C_78_S_4_L_4_out, I5 =>  C_78_S_4_L_5_out, I6 =>  C_78_S_4_L_6_out, I7 =>  C_78_S_4_L_7_out); 

C_78_inst : LUT8 generic map(INIT => "1110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000111010101010100011101010101010001110101010101000") port map( O =>C_78_out, I0 =>  C_78_S_0_out, I1 =>  C_78_S_1_out, I2 =>  C_78_S_2_out, I3 =>  C_78_S_3_out, I4 =>  C_78_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
C_79_S_0_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111011101111111010000000111111111111111011111110111010001111111010000000100010000000000011111111111011101111111010000000111010001000000010000000000000001111111010000000100010000000000010000000000000000000000000000000") port map( O =>C_79_S_0_out, I0 =>  C_79_S_0_L_0_out, I1 =>  C_79_S_0_L_1_out, I2 =>  C_79_S_0_L_2_out, I3 =>  C_79_S_0_L_3_out, I4 =>  C_79_S_0_L_4_out, I5 =>  C_79_S_0_L_5_out, I6 =>  C_79_S_0_L_6_out, I7 =>  C_79_S_0_L_7_out); 
C_79_S_1_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111011101000111111101110100011101010100000001110100010000000100000000000000011111111111111101111111011101000111111101010100011101000100000001110100010000000100000000000000010000000000000000000000000000000") port map( O =>C_79_S_1_out, I0 =>  C_79_S_1_L_0_out, I1 =>  C_79_S_1_L_1_out, I2 =>  C_79_S_1_L_2_out, I3 =>  C_79_S_1_L_3_out, I4 =>  C_79_S_1_L_4_out, I5 =>  C_79_S_1_L_5_out, I6 =>  C_79_S_1_L_6_out, I7 =>  C_79_S_1_L_7_out); 
C_79_S_2_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111111101111111010001000111111111111111011101110100010001111111010001000100010000000000011111111111011101110111010000000111011101000100010000000000000001110111010000000100000000000000010000000000000000000000000000000") port map( O =>C_79_S_2_out, I0 =>  C_79_S_2_L_0_out, I1 =>  C_79_S_2_L_1_out, I2 =>  C_79_S_2_L_2_out, I3 =>  C_79_S_2_L_3_out, I4 =>  C_79_S_2_L_4_out, I5 =>  C_79_S_2_L_5_out, I6 =>  C_79_S_2_L_6_out, I7 =>  C_79_S_2_L_7_out); 
C_79_S_3_inst : LUT8 generic map(INIT => "1111111111111111111111111111111011111111111011101110101010001000111111111111111011101110111010001110100010001000100000000000000011111111111111101110111011101000111010001000100010000000000000001110111010101000100010000000000010000000000000000000000000000000") port map( O =>C_79_S_3_out, I0 =>  C_79_S_3_L_0_out, I1 =>  C_79_S_3_L_1_out, I2 =>  C_79_S_3_L_2_out, I3 =>  C_79_S_3_L_3_out, I4 =>  C_79_S_3_L_4_out, I5 =>  C_79_S_3_L_5_out, I6 =>  C_79_S_3_L_6_out, I7 =>  C_79_S_3_L_7_out); 
C_79_S_4_inst : LUT8 generic map(INIT => "1111111111111111111111111110111011111111111111101110111011101000111111111110111011101110100010001110111011101000100010001000000011111110111011101110100010001000111011101000100010001000000000001110100010001000100000000000000010001000000000000000000000000000") port map( O =>C_79_S_4_out, I0 =>  C_79_S_4_L_0_out, I1 =>  C_79_S_4_L_1_out, I2 =>  C_79_S_4_L_2_out, I3 =>  C_79_S_4_L_3_out, I4 =>  C_79_S_4_L_4_out, I5 =>  C_79_S_4_L_5_out, I6 =>  C_79_S_4_L_6_out, I7 =>  C_79_S_4_L_7_out); 

C_79_inst : LUT8 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000111111101110100011101000100000001111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_79_out, I0 =>  C_79_S_0_out, I1 =>  C_79_S_1_out, I2 =>  C_79_S_2_out, I3 =>  C_79_S_3_out, I4 =>  C_79_S_4_out, I5 => '0' , I6 => '0' , I7 => '0' ); 

 
pred_out <= C_0_out &C_1_out &C_2_out &C_3_out &C_4_out &C_5_out &C_6_out &C_7_out &C_8_out &C_9_out &C_10_out &C_11_out &C_12_out &C_13_out &C_14_out &C_15_out &C_16_out &C_17_out &C_18_out &C_19_out &C_20_out &C_21_out &C_22_out &C_23_out &C_24_out &C_25_out &C_26_out &C_27_out &C_28_out &C_29_out &C_30_out &C_31_out &C_32_out &C_33_out &C_34_out &C_35_out &C_36_out &C_37_out &C_38_out &C_39_out &C_40_out &C_41_out &C_42_out &C_43_out &C_44_out &C_45_out &C_46_out &C_47_out &C_48_out &C_49_out &C_50_out &C_51_out &C_52_out &C_53_out &C_54_out &C_55_out &C_56_out &C_57_out &C_58_out &C_59_out &C_60_out &C_61_out &C_62_out &C_63_out &C_64_out &C_65_out &C_66_out &C_67_out &C_68_out &C_69_out &C_70_out &C_71_out &C_72_out &C_73_out &C_74_out &C_75_out &C_76_out &C_77_out &C_78_out &C_79_out ; 
cor_out <= cor_in; 

end Behavioral;

