--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:25:05 07/27/2019
-- Design Name:   
-- Module Name:   D:/siva/Masters/Thesis/07_ETE_19/part_svhn/svhn_tb.vhd
-- Project Name:  part_svhn
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: SVHN_full_check
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY svhn_tb IS
END svhn_tb;
 
ARCHITECTURE behavior OF svhn_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT SVHN_full_check
    PORT(
         inp_feat : IN  std_logic_vector(511 downto 0);
         out_fin : OUT  std_logic_vector(79 downto 0);
         cor_in : IN  std_logic_vector(79 downto 0);
         cor_out : OUT  std_logic_vector(79 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal inp_feat : std_logic_vector(511 downto 0) := (others => '0');
   signal cor_in : std_logic_vector(79 downto 0) := (others => '0');

 	--Outputs
   signal out_fin : std_logic_vector(79 downto 0);
   signal cor_out : std_logic_vector(79 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: SVHN_full_check PORT MAP (
          inp_feat => inp_feat,
          out_fin => out_fin,
          cor_in => cor_in,
          cor_out => cor_out
        );

   -- Clock process definitions
   --<clock>_process :process
   --begin
		--<clock> <= '0';
		--wait for <clock>_period/2;
		--<clock> <= '1';
		--wait for <clock>_period/2;
   --end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      --wait for <clock>_period*10;
inp_feat <= "11110111111011111111110111110111111011111110111101101011111011101101111101111111111111101101111111111111001101111111111111111101111110111011101100110100110101111111111111011011111011111110110111111111111101011111111111111111110111101010111011011101101011110011111111011111111111111111111011111111101010111111101111111111111111111111110110111110101110111111111001111111101110000110101111110111011101111111111011111111111111111101100111111101101111111111110111111110100111111111111111111111111111001111111111101111";cor_in <= "10110100101101101011101110110111101101100110010010110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11001111111111011111110111011111111111111011111111111111111111111101101111111111011111111111111111111111111101110111011011011111111111111101110111111111111111001111111111110111101111111111010111111111111111110111111111111111111111111101111111111111011111111111101011111101011111011100011111111011011111111111111101111111101110111111111111011111111111111101111111011111110111111111111110111000111111011110111111111111111111110111011111111111011111111101111111111110111111111111111111111101111111111111011111111111";cor_in <= "10110100101101100101111110110111101101101011000110110010101110101011000110110010" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111111111111110111111110110111011011111111111111011111111111101110110111101111111111111111111101111111111111111111111111111010111111011111111111100111110111110111111111001111111101111101111111000111111111111111001001111111111100111111111111111110111111111111111001110101101111111111000101111111011010101111111111101111111110111101111111111111110111111111111111111101111110011111111110111101101111011111111111110111111111111111111011101111111111111111111111110101110111111111111101011111110";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11111111101101111011101011101110111111111111111011111111011101111111000111100100011111111111101111111011111111111011111111111101111101110111111111111111111111111110101111111111011111010101011101110111111111111111111010100111111111111111111110111111111111111001010111110111111110111010111111111111111011001011111111011111000111110110111011111011111011110111110111101111111111111111011111111111111111101110010110111111111011111111101111111011011111111111001100101111111111111110111011011111101111110111011111111110";cor_in <= "01010110101101101011101110110111101101101010010110110010101110101100001010100101" ; wait for 10 ns; 
inp_feat <= "01111110111010101010101111111011100111011110111001101010111101111101011010111101111110111111111111111111101111111011111111111001011011111111111111111001110111111110101110111110001101011111101111010111111011111111111111101111111111111011111111111110111111011111111110011111110110101011111011111111111111011111111111110101111111111111110011110111111111111110110110111111101110001111111111110111111111111011111111111101111110111110110111111111111110011111111111111010110111111111111101111111101111011111111111111011";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111111011111111111111111111111111110111111011111111111110111111111111101011111011111101110110110111111111111111111111111111111111111111111101011111111111111111111111111111101111111111111101111111111111010111100101111111111101110111111101111111101110111111111111111111111111110111111111111111111110111011111110101111110101101011011111111111111111111011110111101111111111111111111111111111110110111111101111111111111101110111111111111111111011101111111111111111111111111111110111111111111011011111010";cor_in <= "11011001101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "01011011111111111111111111111011111110111111111111111111111111111010101111100010111111111111101111101111110111111111111101110111111101111110111010110111111111111111111111111011101111111010001111101110111111111111111111101101111100111111111110111011111111000101101011111111111111111111111011011111111111111111111111111111111111111111111111011010111111111111111011111111111111110110101111111111111101101111111010111111110111111111111111101011101111111111110111101111111111111011111011111111111111110110111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111011101111111110111111110110111111001111111110111011111111110101110110011111111111110110111111111111111111111111101111111011011111111011111011011100111110111110111111111111111101100111101101101111111101111111010101111111111111100111111111111111111111101111111111001110101111111111111010110111011111111111111110001001101101110111101111111111111110011111111111111011111111110010111110101111100100111011111010111110111111111011111111011101111101111110111111111100101011111111111101111011111110";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111101111111111111001011111111111110111111110110111111001110101110111011111111111101110110111111101111111110111111111111110110111111111111111111011111101111110011011100011111111111111111111001111111101111101111111000111110111101010111011111111111101111111111111111111111101111111111001100111101111111111010110111101011110111111111001111101111110111101111111111111110011101111111111011101111111011111111110111101100111010111111111110111111111011111110111101111101011110101111111100101110111111111111001011111110";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11101111111111101100101111111011101011111001111111111111110001000011010110110011111111111111101111011111111111111101111111111101111010110101111011110011111111101110111011110111111111101111101110011101110111111111111111111101111111111111111111111111111111111111110110111111111111111011111111111111011011101111101111111111111111110111111111111111111111111011111101010111111101111111011111111111111111111111111011110011111111010110110101010011110110111101110110110010111111011111110111111111111111111011011111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110100110101110100101" ; wait for 10 ns; 
inp_feat <= "11011111111111011101010111011110011111111011111111111111111110011001110111111110110111111010111011101111011011110111111111101111110110111101111010111101011111111011111111111011111111101100101010111111111111010111111111110110111111101111110011011111111111011111101111111111111111111111111111011011101110111111111111111111111111011111111111111010111011101101111111111111111101110111111111111111111111101111101111111110110111111111011111101011111111011101111111111111111101111111011111111011111111111101111111111111";cor_in <= "10110100101101101011101101011111101101101011000110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "01111110111110101111111111111011101111011111111001111010111101100111011010111001111110111111111111111111111111111011111111111001111011111101111011110101111111111110101111111111011111001111111111010111111111111111111111111111111111111111111111110110011110011011111110111111110111101011111111111111100011111111111011100111111111111111111011111111111111110111110110101111111111111111011111111110111111101111110111111111111110111110110101111111111110001111111110111010110111111111111011111111101111100011111111111010";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11010111111011111110110111110111111111111111111101111011110011001011111111111111111111101110101111111111001001101111111111110101111110111101111111110100100111111111111111111011111011111010110111111111111101111110111011110101111111101011111011010101111011110111111110011111110111111111110011111111101010111111111111111111111111111111110111111110101010101111111111110111111111000110101111111111011101111111111111111111110110111111100111111101111111111111100111110010101111111111111111111110101111010111111111101110";cor_in <= "10110100101101101011101110110111101101100110010010110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111111111111111110111111110111111111001110101110111111111111111101110110011101111111111100101111111101111111111111111111111111011011101011111011011100011011111110111111111101111111111101111111111011111110101111111111001111111111101111101111111111111111101111111111101110111111111110111011111110101011010111111110111111111101110111101101111111111111111011111111111011101101111011111111111111101101111011111011011110111111111111110110001111111101111111110111111101101110111111111111111011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111011111111111111111111111111101011111111111111111111111110111111110110010111011011101010111011111111111111111001111011011111111101010111111111111111010111111111101111111111111011111111111111111111111100101111111111011011111111111011111111111110110111111111011111111111111111111111111111111111111111111101111110111110101110111111111111101010111111111111111111111111011111111111101111101111011111010011101101111101111111101011111111110111100111010111111110001100011111101110111111101111010111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111001111111111111111101111011111011111111111111111111111111111111011111010111001011101010111111111111111111111001111011011111111111010111111111011111110111111111111111111111111011111111111111111011111110101111111111111011111111111011110111111110110111110111011111111111111111111111111101111111101111101011111111111001101110110111111111101010111111011111011101110111011111111111001111101111010111111011111101111101111111111111111111110111101111111111111111101100110110101111111011101111000111011111111011111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111111111111111111111110110111011001111101110111011111111110001110100011111111110101110111011111111111110111011101111111111011111101011111111011100111110111111111111111001111111101111101111111111111110111111011101101111111111100111101111111111111111101111101111011100111111111111111011110111111011110111111110101001101101110111101111111111111110001101111111111111111111111011111111111111100101111011111011111110111111111011111111011101111111001110111111111110111111101111111111101101111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11111110111110101011111110100011101111011110111001111010111001101111011010111101111110111111111111111111111111111011111011111001011111111110111111111101110111111101101110111110011101011111101111010111111111111111111111111111111111111110111111111110011111111011111110011111110111101011111011111110100011111101111011000101111111111101110011110111111111011110110110101101111110011111011111111110111111111011101111111111111110111110110111111101101110101111111111111010110111111111111111111111101111000111111101111011";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111101101011111110111111110111111111111111111111111100110101111111111111110111111111110111111101111010011110101111111111111111111010101111110111101011111111111111111110111111111101101111110111111111110010111011111111111111111101111110011111111111111011111101111111111101111111111111111011011111110110110111000111110111111011101011111101110111111110111101011111111111111111110111111111110111100101111101111111110110101011111011011111101111011111101110111011111111111111111111111011111111111111111111111111111";cor_in <= "10110100101101101011101101011111101101101011000110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111001111111111111111111111111101011110111111111111111111111111111111111111111001111101010111111111111111101111001111011111111111111010111111111111111110111111111111111111111111111111011111111111111111101111111101011111011111111111011111111111110111111111111111111111111111111111111100111110111101111101101111111111011101110111111101111101010111111011111011111110111111111111111101111101111011111011111111111111101111111111111111111111111101111111111111101101100010110101111111111111111111111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111101111111011111110111011111111101100011011111111110111111111101111111111111011111111111110111111101111101111111010010011111101111111111111111111111111111001111111011110111101111111111110111111111111110111111111111011011111110110101111111111011011111111111101011101101011111011111001111111111011101111111011101111011101100111011111111011111111111111100111111011111111111111111101101110000111111111110111101011111101101110111101111111111011111111111111111011111111111111111101111011101111111111111011101111101";cor_in <= "10110100101101100101111110110111101101101011000110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111011101001111110111111101111111011111111011101111111010111110110011111111111111111111001111011111011111111111101111101111111111111111111111111111110101111111111111111110101001101110111111111111111111110110111111111111111110110111101111110111111111111011011110111111000111111111111110011101111011111011111001111111111111111111011111111110110110111101111111111111110111011111111111111111111111110011111111011101111101111111001011111011111001100101111111111111111111111011111101111111111011111101110";cor_in <= "01010110101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111110111111111111111110111111110110111111001110101110111111111111110001110110111101111111111100111111111101110111111111001111111111010110001011110011011100111110111110111111111001111111101111101111111010111110111111010111101111111111101111111111111111110111101111110101011110111111111110110010111111101001110111111110001111111101100111101111111111111111001101111111111010111111110010111111101111101100111011111011111110111111111111111111111101111111111111111111111100101110101111111101101010011111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111101110111111111011111111111111111111111111111111001111111100110111111111111101111101111010111111111111111111111111111111100111010111101111111111111111111111011111011101110111110101011111111110111111111111101111110101111110111111011111111011110101111111111111111111111111111011111001110111111111111111111111111111111101111111010111011111101011111110111111111110110101111111110111101101111111111110111110111111111011111001011111111010111111111111111111111111011111011111101111111111101111111111111";cor_in <= "10110100101101101011101111001111101101101010010110110010101110101011000111010110" ; wait for 10 ns; 
inp_feat <= "10111111111111011101110111011111111011101011011111111111111111111101111111011111011111111111111111011111111101111111010001111111111011111111110111111111111111001110111111111111111111111111110111111111111110111111111111011111111110110101111111111111011111111111001011101001011111011111011111111011011101111111111101111011111110111011111111111111111101111101111111011111110111111111111111111001111111110110111101011111111101111110110111111111111111111111111111111111111111111111111111111111111111111111011101110101";cor_in <= "10110100101101100101111110110111101101101011011110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11010111111011111111110111110101111011111110111101111011111011011111111111110111111111101111110010111111001101111111111111111101111111111010011111110110111111111111111111111111111011111110110111111111111101011111111011111111111111101010111111011101111111110011111111001111111111111111110101111110101010101101101111111111111111111111110110111110101110111111111011111111111110000110101111111111011101111111111111111111110111111111101111101101101111111111110111111010101111111111111111111111111111001110111111101111";cor_in <= "10110100101101101011101110110111101101100110010010111010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111001111111111101111101111011101011110111111111111111011110111101111010011111101111101011111111111011111111111001111011011111111100111111101111111111010111011111111111111111111111111111111111111111111101111110110111111011111111111011111111111110111111111111111111111111111111111111110110110111111111111101111111111011101110111111111111101010111111011111111111111111011111111111001111101111111011111011111101110101111111111111110111111111101111111111111111101100111111100111111111101111111111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111011101111111110111111111110111111001111111110111111111111111101110110111101111111110110111111111111111111111101111111111111011111111011111111011110111111111111111111110001111111101111111111111111111110101111010111101110111111101111101101111111111111111111101111011110101110111111111111111111011011111111111110101001111101100111111111111111111110011111111111111011111111110010111111110111101101111111111011111110111111111011101111011101101111111110111011111100101110111111111111111011101110";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111000011111111111111101111011101011110111111111111111111111111111111011111111001111101010111111111111011011111001111011011111111100011111111111011111110111011110111111111111111111111011111111111111111100101111111111111011111111111011111111111110111111111111111111111111111111111111110111111111101111111101111111111101101110111111111111101010111111011111011111110110011111111111101111101111001111011011111111110101111010101111111111111111101111001111111111101000110110100111111011101111010111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111011011111110111011111111111111111111111111111101111111101111111111111111111111111111111010111101101110111010010111111011111111111111111111111111111001111101111110111111110111111110111111111011110111111111111111111111111110101111111111111011111110111001111110011011111011111001111111111011110111111111101111011101010111110111111011110111111111101111111111111111111111111111110110111111111110110111111111111011001111111111111111110111111111111111111111111111111111111011111111111111111111111111111111111";cor_in <= "11001010101101100101111110110111101101101101100110110010101110101011000110110010" ; wait for 10 ns; 
inp_feat <= "01111110111111111111011111111011111111111111111111111111111101111111110101110010111111111111101011011111111111011111111101111111111110111101101010111111111111101111111111111111101111011111101110001010110111111111110111111101110111111111111110011111011110011111111011111111111111111011111111111111111011111111111111111111111111110111111111011111111111111101011111111111111101110111001111110111111111111111111011111111111111111111110111110011111111111101111111110111111111111111111011111111111111111111111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101110101000101011" ; wait for 10 ns; 
inp_feat <= "11110111101011011111110111011100011111111111101111101111111110011011111111111110110111111110111101101111000011110101111111011111011111011101111110111101111111111011111111111110111011101100101110111111111110110111011111111100111111101111111011111111111011011111111111101111111111111110110111111011101110111110111101111111111111011101111110110110111111111101111111111101111111100100111111111110111100101111101111011110110101111111011111101100011101011101111111111110110101110111011111011011110111011101111111111111";cor_in <= "10110100101101101011101101011111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111110111111111101111111111010101011111101111111011101110101000001011110110011111111111111101111011111111111111011111111111111111010110001111111111111111101111110101111110111111101101111101111011111111011111111111111111101111111111111110111111111111111011011110110111111111111111011111111111111111011101111111111111111111111110111101111111111111110111111111101110111111101011111011111111111111111111111111111111011111111011110110111111111100110011111111110110010111101111111110111111111111111101111011111101111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110100110101110100101" ; wait for 10 ns; 
inp_feat <= "11111110111111101110101111111011101111011110111001111010111011101111011011111101111110111111111111111111111111111011111111111001011011111101111101111100111111111111111110111111011111111111101110000011111111111111111111111111111111111111110111111110110111111011111110011011110111101011111011111110110111111111111111011101111111111101110001010111011111111111110110101111111111011111011111111110111111111011101111111111111110111110111111111111111110001111111100111100111111111111111111111111111111011111111101111110";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111011101101101110111110101111111001111111011101111111011101101101011101111111101111111011110111111111111011111101111101111111111101111111111111111111101111111111001101011111011101110111111111111111111010100110111111111111111110111111111101111101111111111011111100111011111111111111110001111111111101011011100111111110111011011011111111111110110111111111111110111111111111111111111111111111011010011111111011101111101111111011111111111111001101101111111111111111111111011111011101110111111011111110";cor_in <= "01010110101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111111111111111110111111110110111111001110111110111011111111110001010110011101111111110110111111111111111110111111111111111111011111111011110111111100111110111111111111111001111111101111101111111011111110111111111101011111111111101111101111111111111111111111111111001111111111111111111010111111111111010111011110101111101101110111101101111111101110011101111011111111111111111011111111110111101101111011111011111110111011111011111111111111111111011111111111111100101110100111111111101011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11010011111011111111110111110101111111111110111101101011111011011001111101111101111111101111111010111111001101111111111111111101111111111110011111110110111111111111111111011111111011111110110111111111101101011110111011111111111111101011111111010101111011110011111111001111111111011111110101111011101010101101101111111110111111111111110110111110101010111111111011111111111110000110101011111111011101111111111111111111110111111111101011111111101111111111110111111111101111111111111111111111111111001110111111101111";cor_in <= "10110100101101101011101110110111101101100110010010111010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111111111101110111111110110111111001110111110111011111111110101110110111111101110110110111110111111111111111110011111011111011111111011111111011100111110111111111111111001111101101111111111111011111111101111110101001111111111101111101111111111111111101111101111001110111111111111111010111111101011110111111110101111101101100111101111111111111111001111111101111011101111110011111111110111100101111111111011111110111111111111111111011101111111111110111011111110101110111111111101111011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111111111111111111111111110110111111101111111110111111111111110001110110011111111110111110111111011111111111111111111111111111011011111011111110011100111110111110111111111111111111101101101101111111111111111101110101001111111111100111111111111111111111101111111111001110100111111111111011111111111011110101111110011001101101110111101111111111111110101111111111111011111101110011111111101111101101111011111011111110111111111011111111011101111111011110111111111110101110111111111111101011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11101111111111111111110110011111111111110011011111111111111111111001111110111111011111111111110111011111111101111111110111111101111111111111110111111111111110001111111111110111101111111111010111111111111111111111111111101111111110110101111111111111010111111111001011111001011101111111001111111111011101111111011101111111101110111110111111001011111111111110111111011111110111111111111100101100111111010111111101011111111101111110111111111111111111111111011111111111111111111111111111111111111111111111110101111111";cor_in <= "10110100101101100001001110110111101101101010010110110010101110111011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111101111111111011111011111011111111111111111111111011111111110011111111111111101111011111111011011111110101111111111111111111111111110111111111101111111111111111101111111111111110001110111111111111111111101011111101111110111111111111011111011100101011111111111101111011111111011111011111111111111111111111101111110110111111011010111111111111111101011111110111111111101111111111111111011111110011111111111111111110110111111111101111111111111111111110111101111111111111111111111111110101111111111011";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "10111111110111111111101111101111111110111111110110111111001111111110111011111111110101110110011101111111111110111111101101111111111011111111111111011111011011111111011100111101111111111111111011111101101111101101111111111111101111010101001111111111101110101111111111111111111111111111001110101111111111111010111111001011011111111111001001101101110111111011111111111111001001111111111011101111110011111111100111100101111011111111111110111111110010111111011111111111011110101011111100101110111111111111011011111011";cor_in <= "10110100011001101011101110110111101101101010010110111101101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111110111111101110101110111011111011111110111001111010111011101111111110111111111110111111111111111111111111111011111111111001011011111101111011110100111111111111101110110111011010111111101111010111111011111111111111111111111111111010111111111111011111111011111110011101110111101011101011111111110111111111111111111110111011111111110011110111111111111111110110101111101110011111011111111110111111111111111111111111111110110110110111110111111110001111111110111010111111111111111111111111101111101111111101111011";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11011111111111111111111111111111111111011111111111111111111111111011111111101000110111111111101111111111111111111111111101111111011101111110111011110111011111111111111111111111101111111111111111101010111111101111111111101111111110111111111110111011011110011101101111111111111111111111111011011111111111111111111111111111101111111101111111111011101111111101111011111111111011110111101111111111011101111111011111111011111110111110111101101011101111111111111111111111111111111111111111111111111111110111111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "10111111111111011111110110011011111011111111011111111110111111111101111010111111011111111111110111001111111101111111110011111111011111111101110111111111111111001110111111110111101111111111011111111111111111111111111111111111111111110101111111111010001111111111001011111001011111011111011111111111011101111111111101111011111110111110111011011111111111111111111111011111110111111111111110111011111111111110111101111111111101111110111111111111111111111111111111111111111011111111111111111111011111111111111101111101";cor_in <= "10110100101101100101111110110111101101101010010110110010101110111011000110100101" ; wait for 10 ns; 
inp_feat <= "11101110111111111110111111111011111111011111111111111111111101100101011110110011111111111111101111111111111011111011111111111101111011110101111011110011111111111110101111110111111111001111101110010111111111110111111111111111111111111111111111111110011110011011111110111111111111111011111111111111111111011111111111110111111111111111101111110111111111111111110110111111111111111111011111111110111111111111111111111111111111111110110111111111111110001111111110111010111111111111111111111111111111101111011111111011";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111111111111111110111111110110111111001111111110111111111111110001110100011101111111110110111111011111111111111011111111011111011111101011111111011100111111111111111111111001111101111111101101111111111101101111111101101111111111101111111111110111111111111111111111001110101111111111111011110111111011110111111110001011101101110101101111111111111110101101111111111011101111110011111110100111101101111011111011111110111111110111111111011101111111011110111111111100111110111111111101101011101111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "10111111111111011111110111011111111011100011111111111110111111111101111111011111011111111111110111011111111101111111010001111111111111111111110111111111111111001111111011110111101111111111010101111111111100111111111101111011111110110101111111111011001111111111011011100011011111110111001111111011011101111111011101111011101110111111111110011111111101111101111101011111111111111110101111010000111111011110110101111111011011111111111111111111111111111111011111111111111111101111111111101111111111111111011101111110";cor_in <= "10110100101101100101111110110111101101101011000110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "01111111101111111011111011111110111111100111101011101111011101111111010111100010011111111111101111111001111111111011111111111101111101111011111111111111111111111110101111111111011111010001001101010111111111111111111010111111111111111111111110111111111100111001110111110111110110111000111011111111111011001011011111011111100111110111111111111011111011110110110111110111111110011110011111101111111111101111110110111111111011111111101111101010011111111111001101100111111111111111110011011111101101110101011111111110";cor_in <= "01010110101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111110111011101110101110111011111111011110111001111010111011100101111110111101111110111111111111111111111111111011111111111001011011111101111011111101111111111111111011110110011111011111101110000111111111111110111111111111111111111111111111110110010111011011111110011101110111101011111011111111110111111111111111010111111111111101101011110111111111111111110110101111111110011111011111111110111111111111111111111111111110111110111111001111101110101111111110111110110111111111111111111111111111101111111101111010";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11011111111111111111011111011011111111111111111111111111111101011111110111101110111111111111101111101111111111111111111101110111111101111110111010110111111111111111110111111011101111111111001111100110111011111111111111100101111010111110110110110011111111001101101011111101111111111111111111011111111111111111111111111111111111111111111111011011101111111101101111111111111111110110111111111111111111111111111010111111111111111111111111101011101111101111011111111111111101111010111111111101111111110110111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111111111111111111111110110111111001111111110111111111111111100110010011101111110111110111101101101111110110011101111111111011110011011011011111000111111111110111111111001111101111111101101111011111110111011010101001111111111101111101111111111111111111111110111001110101101111111111011111111101001110111111111001101101111110111101111111111111110011101111111111111101111111011111111100111101101111111111111111110111111111111111111101101111111011111111111111110101110110111111111101011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11111111111011111111111111110111111111111110111101111011111011011011111111111101111111101110111010111111001101101111111111111101111110111100001100110100111111111111111111111111111011111110110111111111111101011110111011111111111111101010111011010101111011110111111111001111110111011111110001111111101010101101101111111111111111111111110111111110101100111111111011111101101110001110101111111111011101111111111111111111110111111111101111111101101111111111110111111011101111111111111111111111111111001111111111111111";cor_in <= "10110100101101101011101110110111101101100110010010110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "10111111111101111111111011101111111111111111110110111111001110111110111111111111110101110110011101101111111110111111111111110111111111101111111111011111011011111011011100111110111110111111111101111111101111111111111001101100111111010101101111111111101111111111111111111111101111111111001110101101111111110010111111111111110111111110101111111101100111101111111111111110011101111111111011101111110011111111110111100100111111111011111110111111111011111111011011111111111110100111111100100110111111111101101011111111";cor_in <= "11010010011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11011111111111111101011111111011111111111111111101111111111111011010110111101110111101111111101011110111111111111111111101110111111101111110111010111111111111111111110111111111101011111111101111101010111111111111111111100101110100111110111110111011011111001101111011110111111111111111111101011110111001111111111110111111111110110111111111011011111101111011111011111110111111011111101111110011111111101111111010111011101111111110111111100011101111110111010111101111111111111111111011111111111111110110111111011111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "11111111111011111111110111111101111111111111111111011111111111011001111111111111111111111111111111111111111011111111111111110111111110111100101110111101110101111111111111011011111111111010101111111011110111111111011111111101110110101111111111010111011111010110111011111111111111111111111011111110101111011111111011111111111111111101111111011111101110111101011001111111111111000110111111111111111101111111111111111111111111111111110111101111111111011101111111111110110101111111111111111101111111110111111101111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111011011111111111111111111111111111111111111111101111111111111111111111110111111110111111111111111111111111101011011111111111111111111111111111011110011011110111111111111110111111111111111111111111111111111111111111111111100101111111111111101111111111111111101111111111111111011111111111111111111110110111111111011111111110111111111101110111101111111111111011111011111111111111011111111011110110111111111110101101111011011111111110111111111111111111111111111111111101111111111111111111111101111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000110110010" ; wait for 10 ns; 
inp_feat <= "11111101111011111111110111111111111011111110111101111011111011011011111111111111111011101111111011111111101101111111111111110100111110111100101100110110111111111111111111011011111011111110100111111011111101111111111011111111111111111010111111011111111011110011111111011111110111011111110101111111101010101111101111111110111111111111110110011110101100111111011011111111111110000110101111111111011101111111111111111111110111111111100111111111101111111111110111111010101111111111111111111111101111010111111111101111";cor_in <= "10110100101101101011101110110111101101100110010010111010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10110111111111111011111111111111111111110111111111111111110111111111111111111111111111101111111111111111111101101111111111111111111111111111011111111111111111111111111111111111111111111111110111111111111101111111111111111111111111111111111011011111111111111111111111111111111010111111111111111110111111111111111111111111111111111111111110111111101110111111111111111111101111111111111111110111111111111111111111111111111110111111111111111111110111111111111111111011101011111111111111111111111111010111011110101111";cor_in <= "10110100101101101011101110110111101101101011000110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11111110111111111011110010010111111011110111111111110111111111111101111111110111011111101111111111010111101101111111111011111101111110111111101111111111110111111110111111111111101101111111010111111111111101111111111111101111101110111110111111111111101111110100011011111101010110011111111011111111111111101111111101111111111110111011111110011010101110111111111111011111111111011110111110110011111111111111111010111111111111111111101111111111011111111111111111111111111111111111111111111111111111110111111111110101";cor_in <= "11110000101101100101111110110111101101101100001110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111011111110111010110111111110011011111011111111111111001101111011111011111111011110111111111111111111111010011001111111111111111110111111111110111001111110111111111101111111111010111101111011110111111111111111011111110110101111111111011011111111111001011110001011111110111101111110011011101111111011101111011101100111010011111011011111111011101111111011111111111111111101100110001101111110110111001011111101101111111011111111111111111111111011111111111011011110111111111111111111111111111111101111101";cor_in <= "10110100101101100101111110110111101101101011000110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111111011111111111111111111111111111101111010111111100010111111111111101111001111111111111111111101110111111101111010111110110111111111111111111111111111101111111011011111001010111111111111111011100101111110111111111110111111011111011101101011111111111101111111111011011110111011111111111111111101101111110111111111011011101001111111111001111110111111010111101111110111011111101111111010111011111111111110111111100011101111011101111111111111110101111111111001111111111110110111111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "10011111111111011110110111010111111011111011011111111110111111111001100011111111011111111011110111011111111101111111010011101111011111111111110111111111111111001110111111110111101111111111111111111111111110111111111111111111111110110101111111111011011111111111101011111001011111011011011111111111011101111111111101111011101100111011111111011110111110011101111111011111111111111111111110110001111111011110111001011111111101111111111111111111111111111011111111111111111011111111111111111101111111111111111101111101";cor_in <= "10110100101101100101111110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111011111111111101111101111111101011110111111111110111111110111111011111011111001011101010111111111111111111111001111011011111111101011111111111011011010111111111101111110111111111111111111111111111011101101111111111111011111011111011111111111110111111111111111111111111111111111111110111111111101111111111111110111111101111110111101111101010111111011111110111011111011111111111001111111111111111111011111111101101111111111111111111111110101111111111111111001100011111101111111111111111110111111011111111011";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111101111111111011111111011111101111110110111111001111111110111111111111111001110110011101111111110110111111111111110111111111111111111111011111111011110011011100111111111111111111111001111111101111111101111111101110111001110111101111111111101111101111111111111111101110101111001110101111111111111011110111101011110111111110001111101101110111111111111111111100001111111111110011101111111010111111101111101101111011111011111110111111111011111111111001111111011110111111111100101110111111111111101011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11011111100111111111011111111110111111111111101111101111111111111111001111100110010111111111111111110111111011111111111111111101111111111111111011111111111111111111111111011111111101110101001100110111111111111111111111110111111111101111111111110111111111011101111111110011111111111011111111111111101111011111111101111111101111111110111010111011111011110101110111111111111111111111111111111111111111101111010110111111111111111111101111101010011111011111011111101111111101111111111011011111101101110111111110111110";cor_in <= "01010110101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111110101101101111101111111011111111011110101111111010111111100111011110111111111110111111111111111111111111111011111111111101011111111111111111111101111111111111111111111111011111001111101100010111111111111111011111111111111111111111111111111110110111011111111110111111110111101011111111111110111111011111111111010111111111011111110111111111111111111111110110111111111111011111011111111110111111111111111111111111111010111110111111011111111110001111111111111110111111111111011101111111111111011111111111111110";cor_in <= "10110100101101101011101111001111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11010011111111111101111111011011111111110011111111111111111101011011100111100010111111111111101111001111111111011111110101110111111101110110111010110111111111111111111111111111101011111011001111101010110111111111111111101101111110111110111110111011111111001101101011111111111111111111111111011111111011111111111111111111111110110111111111011010001011111101011001111111111111110110101111111011111111101111011010111111101111111111111111101011101111111111110111111111111101111111111011111101111111110110111111111101";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000101101100" ; wait for 10 ns; 
inp_feat <= "11011111101111011101110111111100011101111011011111111111101110010101111111111111110111111111111011101111010011110101111111111111110111010101111111111111111111111011111111110111111011101100101110111111111111011111011111010110111111101111110011111111011011010111101111111111011111110111110111011011111111110110111001111111011111011101111110111110111111111111101111111111111111100100111001111111111100101111101111011110110101011111011111001100011111111101111111111111110110111111011111011011111111111101111111111111";cor_in <= "10110100101101101011101101011111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111011111110110011111111111111011011111111111111111111101111111111111011111111111110111111111111001110111011011011111111111111101110111111111111111001111111111110111101111111111110010111111111110111110111111111011111110110101111111111111001111111111111011101001011111011111001111111011011101111111111001111011111110111110111111011111111111101101111111011111110111110111111110010001111111111110111101011111111101111111011011111110111111111101111111111111111101111111111111111100111111111111111101111101";cor_in <= "10110100101101100101111110110111101101101010010110110010101110111011000110100101" ; wait for 10 ns; 
inp_feat <= "11011111111111011110110111011101011101111111111111111111110110111111111111101111111111111111111101101111111111110111111111100111111110110101111110111101111010110011111101111111111111101110101010111111011111111111111111110100111111101111111011011111111111111111101111111111111111110111110111111111101110111111111111111111111111011111111111111110111011101111111111111101111101100111111111111111111111101111111110111110110101111101011111101110111111011101111111111111111111110111011111111011111011111101111111111111";cor_in <= "10110100101101101011101101011111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11110111011011111101110111110111111111111110111111111010111011011001111111111101111111101111111011111111001001111111111111111001111111111101011101110110111111111111110111111011111011111110110111111111111101011110111111111111111111101011111011110101111011110011111110001111111101011111110011110111101110101111101111111111111111111111110110111110101110101111111101111101111110000110101011111111011101111111111111111111110111111111100111111101101111111110111111111011101111111111111111111111111111001111111111111111";cor_in <= "10110100101101101011101110110111101101100110010010111101101110101011000110110010" ; wait for 10 ns; 
inp_feat <= "11111111111111111111011011101111111111101111110010111111001111111110111111011111111010110110011111111111111110111111011111110111111011111111011111011111111111111111111100111111111111111111111101101111111111101111111111101111111011111101101110111111100111101111111111111111101111111111001110111101111111111011110111101011010111111110001101111101110111111111111111101110001101111111111011101111110010111110111111100111101010111011111110111011111011111110111111111101011010101011111110100110111111111111101011111011";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111111111111111110111111110110111011001111101110111111111111110111110110011100111110101110111111011111111110111111111111111111011011001011011011011000111110111110111111111001111101101111101101111110111110101111110101001111111111101111101111111111111111111111111101001110111111111110111010111111111011110101111110101111101111110111101111111111111110101101111111111011101111110010111111111111101100111011111011111110111111111011111111001101111111111110111111111100101110111111111111101111111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111011011111111111111100111111101011110111111111110111111111111111111111011111011101101010111111111011011111111001111011011111111111000111111111111111010111111111111111111101111111111111111111111111111100101111111111111011111111111011111111011110110111110111011111111111111111110111110111111111111111101101111111111001101010111111111111101011101111011111011111111111011111111101101111101111101101011011111111111101111111111111111111110111100111011111111111001100111111101111111111101111010111011111111011111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111110111011101110101111111011111011011110111001111000111011100101011011111101111110111111111111111111101111111011111111111001011011101111111111110101110111111111101011111101001011110111111111000111111011111111111111111111111111111010111111111110111111111011111110011111110111101011111011111110100011011111111111110101111011111111100011110111111111111011110110111111111111011111011111111110111111111111111111111111111110111110110111111111101110000111111110111010110111111111111101111111101111001111111101111011";cor_in <= "10110100101101101011101110110111101101101010010101101110101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10001111111011011111110111011111111011111011111111111111111111111001111111111111010111111111110111011111111101111111010001111111111111111111111111110111111111001111111111110111101111111111110111111111111110111111111111111011111110110101111111111111001111110111001011111101011111010111001111110011011101111111111101111011101110111011111110011111111110101101111111011111111101111111111110110111111111110110111011111011111101111111011011110111111111110111111111111111111101111111011111111111111111111111111101111101";cor_in <= "10110100101101100101111110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111110111111111011111011111101111111101101110101111111111010110011101111111111101111011111111111111111111111111101111110110011101011111111110111111111101111111111101101011111111111011111111011111111111111101101111111111111111111111111011110011111111010111111111110111011111111111111110111001111111111110111111111110111111111010111111110111111111101010111111111111111111111110111111111111111111011111111111111111110100111111111100111111111111111110010110111111111110101111111111111110111011111111011";cor_in <= "10110100101101101011101110110111101101101010010110110010101110100110101110100101" ; wait for 10 ns; 
inp_feat <= "11010111101111011101110111111101011111111011111111111111100110011001111111111110110111111110111101101110010011110101111111011111111111110101111010111101101111111011111111111111111011101110101010111111111111010111011111110101111111101111110011111101011111011111101111101111111111110111110111011011101110111111111111111111111111011101111111111110111111111111001011111111111111100110111111111111111101100111101111111110111111111111011111001100111011011101111111111111110101111111011111111011111011111101111111111101";cor_in <= "10110100101101101011101101011111101101101010010110110010101110111011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111011101111111110101111110010111111001111111110110111111111110001110100011100111111111110111111011111111110111111111111111111011110011011111111011100111110111111111111111101111011101111101111111101111111101111110111001111111111101111101111111111111111101111111111001100101111111111111010110111111011110111111110001001111101110111111111111111101110011111111111110111111101111011111111111111100101111011111011111110111111111011111111001101111111111110110111111100101111110111111111101011111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11111111011111111111101111101111111101011110111111111111111111110111111010110111111001011101010111111011111111111111001111011011111111101011111111111111111110111111111111111101111111111111011111111111111111100101111111011111011111111111011111111111110111111111111111110111111111111111111111111111111111111101101111110111001101110111111101111101010111111111111111111101111011111111011101111101111001111111011111101111101111111111111111111111111100111011111111111101100110110100111111011111111010111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111101111111110111111111110111011001110111110111111111111110100111110111111111011111111111111111111111111111111111111111111011111111011111011101100111111011111111110111101111111111111111101111011111110111111111111101111111111101110111111110111111111110111111111111111111111111111111011111111011111111111111111111111111101110111101111111111111110001010111011111011101111110111111111111111111101111111111011111110111011110111111110001101111111111111111111111101101111111111111111111111111110";cor_in <= "10110100011001101011101110110111101101101010010110111101101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "10110101111100111011111011110110111111101111011111101111110111111111101110011111101111111111011111111111110111110101110111110111111111111111000110111101111111111111110111111110111111111111111111111110011110111111111111111111110011110111101011011110111111111111001111111111111110110111110111101111111111110111111111111110110110111011011111111111111111011111111111111101101111111111111110110111101111111111001001011011111101111101111111110111011111111111111111101111111011111111111111110111110011011111101011001101";cor_in <= "10110100101101101011101110110111101101101010010110110010011010001011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111111111111111111111111111111101111111110111111001111111110111111111111110011010110011101111111110110111111111111111111111111111111111111011111011111110011111111111111111111111111111111111110101111111111111011101100111101110111101111111111111111111111111111111111111110110111111111111111111111110110111111111111111101111110001101111111111111101111111110111110011111111111111011111111111110111111111111111111111101111011111110111111111011110111001111111111111111111111111101111110111111111111101111111111";cor_in <= "10110100011001101011101110110111101101101010010110110010111001001011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111011101110110011111111011111011111111111111111111111111111101010111011111111111110111011101111101110111010001011111111111111111110111111111111111001110111011110111111110111111111111111111111110111111111111011111101101110101111111111111011111111111101011111001011111011111011111111011011101111111111111111011101110111110111111011111111111111111111111011111111101111111111110110101101111110110111101011111101101110111111111110111111111111011111111111111111111111111111111011111111111111111011111111101";cor_in <= "10110100101101100101111110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111101111111111111101101111110111111110110111111001111101110111111111111110101010110011101111110110110111111111111111111111111111111111111011110011011111011011100111110111111111111111001111111101111101101111100101111111111111111001111111111101111101111111111111111101111111111001100101111111111110000111111101011110111111110101111101101110111101110111111101110001111111111111111101111111011111011100111100100111011111011111110111111111111111110111111111101011110111111111100101110111111111111111011011111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11110110111101111011111010110110001111110111011111101111110111111111111110011111101010111111111111111111110111110101100111111111111111111111010110111101111111111101110111111110111111111111111111111010011110111101111111101111110010111111111011011110111111111110111111111111110100110111110111101101111111010111111111011111111110111011011111111111111111111111111111111101100111111111111111100111101111111111101101011011111111111111111111110111100111111111110111101011111011110111111111111111110011011111101111011101";cor_in <= "10110100101101101011101110110111101101101010010110110010011010001011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111110111111111111011111111111110101111110010111111001111111110111111111111110001010110011101111110110110111111111101111110111111111111111111011111011011110111011100111010011111111111111101111111101111101111111010111110111111111111101111111111100111100101110111111111101111111111111100101111111111111000110111111001010111111111101001101111110111101111111111101110001100111111111011101111111011111110110111101101111010111011111110111111111111111110001101111101011110111111111100101110111111111111001011001110";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "01111111111111111011101010111110111101110111111011101111011111111111010111110110111111111111111111111001110111110111111111111101111101111011111101111111111111111111111111111111111111110101001101110111111111111111111111110110111111111110111110111111111111111101111111110011111110111110111011111110111011101111011111011111100111111110111110110011111011110111110111110110111111111111111111111111011111101111011110011111111111111111101111101011011111111010001101101110111111111100111111011111101111110011111111101110";cor_in <= "01010110101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111111011111111011111111111110110111111101111111110111110111111111101111110011111111111111100111111111011111110111011111111111111011011011011011111011110111110111111111111111011111111101111111111111110111111101111110101101111111111111111111111111111111111111111111111001110111111111111111011110111111011110111111110001011111101110111111111111111101111001111111111111011111111110011111110101111100110111010111011111111111111111011111111011111111111111110111111111100111111111111111111001111111111";cor_in <= "10110100011001101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11110111010111111111111111101111111101011110111111010111111111111111101011111010111011011101010101111111111111011111001111011111111111101010111111111111111010110011110101111111101111111111111111111111111111100101111111111111011111111111111111101111110111111111111111110111111111111111111110011111111111111111111111110111000101110111011101111101011111111111111111111110110011111111111101111101111011111011011111101111101111111111011110111111111101111011111111111101100111110101111111111111111010111111111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111011111111111111111100111011101011110111111011111111011111111111111111111111101111101010111111101111011111111001111011011111111101010111111111111111110111111111111111111111111111111011111111111111101100111111110111111011111111111011111111011110111111111111011111110111111111111111101011111111101111111101111111111101101110101111101111101011111111111111011111111111011110111101101111101011010111111011111111111101111111111011111111111111101111101111111111001100011110101111111011101111010111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111110111011111111111111111111101111111110111101111001111011111101111110111111111111101111111111111111101111111011111111111001111111111110011101111110111111111111111111111111111011111111111111011111111111111111111111111111111111111111111111111101111111110111111111011111110111111011111111111111111011111101111111111110111111111011110111111111111110111111111111111111111110011110011111111111111111111111111111110111111110111110111111111111101110101111111111111110111111111111111111111111011111001111111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111001110111111111111101111111101011110111111111110111011110111111011101010111001111101010111111111111111111111001111011011111111110010111101111111110110111111110111111111111111111111011111111111111101100101111110111111011111111111011110111010110111111111111011111111111111111111111110011110101101111111001110110111001001110111111101111101010111111011111010111110111011110111111101111101111011111011011111111111101111111101111111111110111101111011111111111101100110110101111111111101111010111011111111111111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111011111111111111111101111111101011110110111111111111011111111111011111110111001101101010111111011111111111111001111011011110111111010111111111111111010111111111101111111111101111111011111111111111111100101111110111111011111111111011111111111110110111111111011111111111111111111111110001111111111111111101111110111010101110110111111111101010111111011111011101110111011111111111101111101111011111011011111101111101111111111111111111110111101111010111111111001100010110101111111111101111010111011111111110111";cor_in <= "10110100101101101011101110110111011011001010010110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "10111111111111111111110111010111111011111001010111011110111111111101111111011111011101111111110111111111111101110111011011111111111111111111111111111111111111001111111011110111111111111111110111111111011110101111111111011111111100110101111111111011011111111111101011101001011111011101001111111011011101111111011111111011101110111111111111011111111101011101111111011111111101111101111101111001111111010100111101111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111101111101";cor_in <= "10110100110010010101111110110111101101101011000110110010101110101011000110100101" ; wait for 10 ns; 
inp_feat <= "11110111111101111111111111111010111111111111111111101101100111111111101010110111101111111111111111011111111111110111101111111111111111111111010111111111111111111111111111111111101111011111111111111111011110110111111111101111110111111111111111111110111111111111111111111111111110110111111111111111111111011111111111111111111111111111011111111111111111111111111111111111111101111111011111100111111111111111111101111011111111011111111110110111111111111111111111111011111011111101111111111111110011111111111111111111";cor_in <= "10110100101101101011101110110111101101101010010110110010111000011011000110100101" ; wait for 10 ns; 
inp_feat <= "11111111111101111111111111101111101111111111110110111011001111111110111111111111110001110110011100111111110110111111011111111110111111111111111111011111111011111111011110111111111111111111111101111101101111101111111110111111111111011111011111111111100111101111111110111110101111101101101100101111111111111100111111111011011111111111001001111101110111111111111111111110001111111111111011111111111010111111110111101101111110111011111100111111111010111111111101111111111110111111111110101111101111111111101011111010";cor_in <= "10110100011001101011101110110111101101101011000110110010101110101011000110110001" ; wait for 10 ns; 
inp_feat <= "11110111111101111011111111110110111111111111011111111111110111111111101110011111101110111111111111011011111111110111110111111111111111110111000111111111111111111101110111111110111111111111101111111110011110111101111111111011110011111101111011011111111101111111011111111111111000110111110111111111111111000111111111111111111110111011011111111110111110111111111111101101101111111111111111000111101111111111001101011011111101011111111011110111100111111111111111101111111011111111111110111111110010011111101111011101";cor_in <= "10110100101101101011101110110111101101101010010110110010011010001011000110100101" ; wait for 10 ns; 
inp_feat <= "10110101111101111011111011110110111111100011011111011111110111111111111110011111101110111111011111111111111111110111110111111111111111111111010110111111111111111111110111111110111111111111111111111110011110111101101111111111110011110101111011011111111111111111001111111011011000110111110111111011111111010111111111111110110110111011011111111110111111011111111111111101101111111111111110000111101111111011101101011011111100111111111111110111101111111101111111101111111011110111111110111111110010011111101111011101";cor_in <= "10110100101101101011101110110111101101101010010110110010011010001011000110100101" ; wait for 10 ns; 

      -- insert stimulus here 

      wait;
   end process;

END;
