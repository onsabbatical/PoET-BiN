----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:12:42 07/23/2019 
-- Design Name: 
-- Module Name:    cifar_fin_layer - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cifar_fin_layer is
    Port ( inp_feat : in  STD_LOGIC_VECTOR (79 downto 0);
           cor_in : in  STD_LOGIC_VECTOR (79 downto 0);
           cor_out : out  STD_LOGIC_VECTOR (79 downto 0);
           out_fin : out  STD_LOGIC_VECTOR (79 downto 0));
end cifar_fin_layer;

architecture Behavioral of cifar_fin_layer is
component LUT8
generic(INIT : std_logic_vector(255 downto 0) := (others => '0') );
port(I0:in std_logic;
I1:in std_logic;
I2:in std_logic;
I3:in std_logic;
I4:in std_logic;
I5:in std_logic;
I6:in std_logic;
I7:in std_logic;
O:out std_logic);
--  Port ( );
end component;

signal C_0_B_7_out : std_logic := '0'; 
 signal C_0_B_6_out : std_logic := '0'; 
 signal C_0_B_5_out : std_logic := '0'; 
 signal C_0_B_4_out : std_logic := '0'; 
 signal C_0_B_3_out : std_logic := '0'; 
 signal C_0_B_2_out : std_logic := '0'; 
 signal C_0_B_1_out : std_logic := '0'; 
 signal C_0_B_0_out : std_logic := '0'; 
 signal C_1_B_7_out : std_logic := '0'; 
 signal C_1_B_6_out : std_logic := '0'; 
 signal C_1_B_5_out : std_logic := '0'; 
 signal C_1_B_4_out : std_logic := '0'; 
 signal C_1_B_3_out : std_logic := '0'; 
 signal C_1_B_2_out : std_logic := '0'; 
 signal C_1_B_1_out : std_logic := '0'; 
 signal C_1_B_0_out : std_logic := '0'; 
 signal C_2_B_7_out : std_logic := '0'; 
 signal C_2_B_6_out : std_logic := '0'; 
 signal C_2_B_5_out : std_logic := '0'; 
 signal C_2_B_4_out : std_logic := '0'; 
 signal C_2_B_3_out : std_logic := '0'; 
 signal C_2_B_2_out : std_logic := '0'; 
 signal C_2_B_1_out : std_logic := '0'; 
 signal C_2_B_0_out : std_logic := '0'; 
 signal C_3_B_7_out : std_logic := '0'; 
 signal C_3_B_6_out : std_logic := '0'; 
 signal C_3_B_5_out : std_logic := '0'; 
 signal C_3_B_4_out : std_logic := '0'; 
 signal C_3_B_3_out : std_logic := '0'; 
 signal C_3_B_2_out : std_logic := '0'; 
 signal C_3_B_1_out : std_logic := '0'; 
 signal C_3_B_0_out : std_logic := '0'; 
 signal C_4_B_7_out : std_logic := '0'; 
 signal C_4_B_6_out : std_logic := '0'; 
 signal C_4_B_5_out : std_logic := '0'; 
 signal C_4_B_4_out : std_logic := '0'; 
 signal C_4_B_3_out : std_logic := '0'; 
 signal C_4_B_2_out : std_logic := '0'; 
 signal C_4_B_1_out : std_logic := '0'; 
 signal C_4_B_0_out : std_logic := '0'; 
 signal C_5_B_7_out : std_logic := '0'; 
 signal C_5_B_6_out : std_logic := '0'; 
 signal C_5_B_5_out : std_logic := '0'; 
 signal C_5_B_4_out : std_logic := '0'; 
 signal C_5_B_3_out : std_logic := '0'; 
 signal C_5_B_2_out : std_logic := '0'; 
 signal C_5_B_1_out : std_logic := '0'; 
 signal C_5_B_0_out : std_logic := '0'; 
 signal C_6_B_7_out : std_logic := '0'; 
 signal C_6_B_6_out : std_logic := '0'; 
 signal C_6_B_5_out : std_logic := '0'; 
 signal C_6_B_4_out : std_logic := '0'; 
 signal C_6_B_3_out : std_logic := '0'; 
 signal C_6_B_2_out : std_logic := '0'; 
 signal C_6_B_1_out : std_logic := '0'; 
 signal C_6_B_0_out : std_logic := '0'; 
 signal C_7_B_7_out : std_logic := '0'; 
 signal C_7_B_6_out : std_logic := '0'; 
 signal C_7_B_5_out : std_logic := '0'; 
 signal C_7_B_4_out : std_logic := '0'; 
 signal C_7_B_3_out : std_logic := '0'; 
 signal C_7_B_2_out : std_logic := '0'; 
 signal C_7_B_1_out : std_logic := '0'; 
 signal C_7_B_0_out : std_logic := '0'; 
 signal C_8_B_7_out : std_logic := '0'; 
 signal C_8_B_6_out : std_logic := '0'; 
 signal C_8_B_5_out : std_logic := '0'; 
 signal C_8_B_4_out : std_logic := '0'; 
 signal C_8_B_3_out : std_logic := '0'; 
 signal C_8_B_2_out : std_logic := '0'; 
 signal C_8_B_1_out : std_logic := '0'; 
 signal C_8_B_0_out : std_logic := '0'; 
 signal C_9_B_7_out : std_logic := '0'; 
 signal C_9_B_6_out : std_logic := '0'; 
 signal C_9_B_5_out : std_logic := '0'; 
 signal C_9_B_4_out : std_logic := '0'; 
 signal C_9_B_3_out : std_logic := '0'; 
 signal C_9_B_2_out : std_logic := '0'; 
 signal C_9_B_1_out : std_logic := '0'; 
 signal C_9_B_0_out : std_logic := '0'; 
 
 
 signal C_0_out : std_logic := '0'; 
 signal C_1_out : std_logic := '0'; 
 signal C_2_out : std_logic := '0'; 
 signal C_3_out : std_logic := '0'; 
 signal C_4_out : std_logic := '0'; 
 signal C_5_out : std_logic := '0'; 
 signal C_6_out : std_logic := '0'; 
 signal C_7_out : std_logic := '0'; 
 signal C_8_out : std_logic := '0'; 
 signal C_9_out : std_logic := '0'; 
 signal C_10_out : std_logic := '0'; 
 signal C_11_out : std_logic := '0'; 
 signal C_12_out : std_logic := '0'; 
 signal C_13_out : std_logic := '0'; 
 signal C_14_out : std_logic := '0'; 
 signal C_15_out : std_logic := '0'; 
 signal C_16_out : std_logic := '0'; 
 signal C_17_out : std_logic := '0'; 
 signal C_18_out : std_logic := '0'; 
 signal C_19_out : std_logic := '0'; 
 signal C_20_out : std_logic := '0'; 
 signal C_21_out : std_logic := '0'; 
 signal C_22_out : std_logic := '0'; 
 signal C_23_out : std_logic := '0'; 
 signal C_24_out : std_logic := '0'; 
 signal C_25_out : std_logic := '0'; 
 signal C_26_out : std_logic := '0'; 
 signal C_27_out : std_logic := '0'; 
 signal C_28_out : std_logic := '0'; 
 signal C_29_out : std_logic := '0'; 
 signal C_30_out : std_logic := '0'; 
 signal C_31_out : std_logic := '0'; 
 signal C_32_out : std_logic := '0'; 
 signal C_33_out : std_logic := '0'; 
 signal C_34_out : std_logic := '0'; 
 signal C_35_out : std_logic := '0'; 
 signal C_36_out : std_logic := '0'; 
 signal C_37_out : std_logic := '0'; 
 signal C_38_out : std_logic := '0'; 
 signal C_39_out : std_logic := '0'; 
 signal C_40_out : std_logic := '0'; 
 signal C_41_out : std_logic := '0'; 
 signal C_42_out : std_logic := '0'; 
 signal C_43_out : std_logic := '0'; 
 signal C_44_out : std_logic := '0'; 
 signal C_45_out : std_logic := '0'; 
 signal C_46_out : std_logic := '0'; 
 signal C_47_out : std_logic := '0'; 
 signal C_48_out : std_logic := '0'; 
 signal C_49_out : std_logic := '0'; 
 signal C_50_out : std_logic := '0'; 
 signal C_51_out : std_logic := '0'; 
 signal C_52_out : std_logic := '0'; 
 signal C_53_out : std_logic := '0'; 
 signal C_54_out : std_logic := '0'; 
 signal C_55_out : std_logic := '0'; 
 signal C_56_out : std_logic := '0'; 
 signal C_57_out : std_logic := '0'; 
 signal C_58_out : std_logic := '0'; 
 signal C_59_out : std_logic := '0'; 
 signal C_60_out : std_logic := '0'; 
 signal C_61_out : std_logic := '0'; 
 signal C_62_out : std_logic := '0'; 
 signal C_63_out : std_logic := '0'; 
 signal C_64_out : std_logic := '0'; 
 signal C_65_out : std_logic := '0'; 
 signal C_66_out : std_logic := '0'; 
 signal C_67_out : std_logic := '0'; 
 signal C_68_out : std_logic := '0'; 
 signal C_69_out : std_logic := '0'; 
 signal C_70_out : std_logic := '0'; 
 signal C_71_out : std_logic := '0'; 
 signal C_72_out : std_logic := '0'; 
 signal C_73_out : std_logic := '0'; 
 signal C_74_out : std_logic := '0'; 
 signal C_75_out : std_logic := '0'; 
 signal C_76_out : std_logic := '0'; 
 signal C_77_out : std_logic := '0'; 
 signal C_78_out : std_logic := '0'; 
 signal C_79_out : std_logic := '0'; 
begin

C_0_out <= inp_feat(0); 
C_1_out <= inp_feat(1); 
C_2_out <= inp_feat(2); 
C_3_out <= inp_feat(3); 
C_4_out <= inp_feat(4); 
C_5_out <= inp_feat(5); 
C_6_out <= inp_feat(6); 
C_7_out <= inp_feat(7); 
C_8_out <= inp_feat(8); 
C_9_out <= inp_feat(9); 
C_10_out <= inp_feat(10); 
C_11_out <= inp_feat(11); 
C_12_out <= inp_feat(12); 
C_13_out <= inp_feat(13); 
C_14_out <= inp_feat(14); 
C_15_out <= inp_feat(15); 
C_16_out <= inp_feat(16); 
C_17_out <= inp_feat(17); 
C_18_out <= inp_feat(18); 
C_19_out <= inp_feat(19); 
C_20_out <= inp_feat(20); 
C_21_out <= inp_feat(21); 
C_22_out <= inp_feat(22); 
C_23_out <= inp_feat(23); 
C_24_out <= inp_feat(24); 
C_25_out <= inp_feat(25); 
C_26_out <= inp_feat(26); 
C_27_out <= inp_feat(27); 
C_28_out <= inp_feat(28); 
C_29_out <= inp_feat(29); 
C_30_out <= inp_feat(30); 
C_31_out <= inp_feat(31); 
C_32_out <= inp_feat(32); 
C_33_out <= inp_feat(33); 
C_34_out <= inp_feat(34); 
C_35_out <= inp_feat(35); 
C_36_out <= inp_feat(36); 
C_37_out <= inp_feat(37); 
C_38_out <= inp_feat(38); 
C_39_out <= inp_feat(39); 
C_40_out <= inp_feat(40); 
C_41_out <= inp_feat(41); 
C_42_out <= inp_feat(42); 
C_43_out <= inp_feat(43); 
C_44_out <= inp_feat(44); 
C_45_out <= inp_feat(45); 
C_46_out <= inp_feat(46); 
C_47_out <= inp_feat(47); 
C_48_out <= inp_feat(48); 
C_49_out <= inp_feat(49); 
C_50_out <= inp_feat(50); 
C_51_out <= inp_feat(51); 
C_52_out <= inp_feat(52); 
C_53_out <= inp_feat(53); 
C_54_out <= inp_feat(54); 
C_55_out <= inp_feat(55); 
C_56_out <= inp_feat(56); 
C_57_out <= inp_feat(57); 
C_58_out <= inp_feat(58); 
C_59_out <= inp_feat(59); 
C_60_out <= inp_feat(60); 
C_61_out <= inp_feat(61); 
C_62_out <= inp_feat(62); 
C_63_out <= inp_feat(63); 
C_64_out <= inp_feat(64); 
C_65_out <= inp_feat(65); 
C_66_out <= inp_feat(66); 
C_67_out <= inp_feat(67); 
C_68_out <= inp_feat(68); 
C_69_out <= inp_feat(69); 
C_70_out <= inp_feat(70); 
C_71_out <= inp_feat(71); 
C_72_out <= inp_feat(72); 
C_73_out <= inp_feat(73); 
C_74_out <= inp_feat(74); 
C_75_out <= inp_feat(75); 
C_76_out <= inp_feat(76); 
C_77_out <= inp_feat(77); 
C_78_out <= inp_feat(78); 
C_79_out <= inp_feat(79); 


C_0_B_0_inst : LUT8 generic map(INIT => "0100110010011001011011001101100110110011011001101001001100100110110011011001100101001100100110010011001001100110101100110110011000110110011001000011001001100110110010011001101111001101100110010010011001101100001101100110010011011001100100111100100110011011") port map( O =>C_0_B_0_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_1_inst : LUT8 generic map(INIT => "1000000000010001011111111110111000110011011101111110110011001000111111101110111010000000000100011100110010001000001100110111011100110111011101111100110010001000111111101110110000000001000100011100100010000000001101110111011100010001000100111111111011101100") port map( O =>C_0_B_1_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_2_inst : LUT8 generic map(INIT => "1100001100101101101111001100001100001111101101001100001100111100001111001100001100111100110100101100001100111100111100000100101100001011101101001100001100111100001111001100001100111101110100101100001100111100111101000100101100101101110100001100001100111100") port map( O =>C_0_B_2_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_3_inst : LUT8 generic map(INIT => "1100000011111101000000111100000011111111000010111100000011111100111111000011111100000011110100000011111100000011111100001011111100000000111101000011111100000011111111000011111100000010110100001100000011111100000010110100000011111101001011111100000011111100") port map( O =>C_0_B_3_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_4_inst : LUT8 generic map(INIT => "0110101001010111101010100110101010101010101010101001010110101001101010011010101001010101100001010101010101010101010110100101010101010101101000010101010101010101010101100101010110101010011110100110101001010110101010101110101010101000101010101001010110101001") port map( O =>C_0_B_4_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_5_inst : LUT8 generic map(INIT => "0001101000001111010110100001101001011010010110100111000001011000101001111010010100001111100011110000111100001111000010100000111100001111101011110000111100001111000011100000111101011010000010101110010111110001101001011110010110100111101001011000111110100111") port map( O =>C_0_B_5_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_6_inst : LUT8 generic map(INIT => "0000101000001111000010100000101000001010000010100000000000001000101011111010111100001111100011110000111100001111000010100000111100001111101011110000111100001111000011100000111100001010000010101110111111111111101011111110111110101111101011111000111110101111") port map( O =>C_0_B_6_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 
C_0_B_7_inst : LUT8 generic map(INIT => "0000101000001111000010100000101000001010000010100000000000001000101011111010111100001111100011110000111100001111000010100000111100001111101011110000111100001111000011100000111100001010000010101110111111111111101011111110111110101111101011111000111110101111") port map( O =>C_0_B_7_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out, I6 =>  C_6_out, I7 =>  C_7_out); 

C_1_B_0_inst : LUT8 generic map(INIT => "0000010110101010101010100101111101011111101001011010010101011010010111111010010110100101010110100101101000000101000001011010000000000101101010101010101001011111010110101010010110100101111110100101111110100101101001010101101001011010010101010000010110100000") port map( O =>C_1_B_0_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_1_inst : LUT8 generic map(INIT => "0011110001101001100101100011110011000011100111000110001111000110001111000110001110011100001110011100011000111100110000111001110000111100011010011001011000111100110001101001110001100011110001100011110001100011100111000011100111000110001111001100001110011100") port map( O =>C_1_B_1_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_2_inst : LUT8 generic map(INIT => "1001010110000001111010000110101001010110000101011000100110101000011010100111011000010101100100011010100001101010010101100001010110010101100000011110100001101010010101110001010110001001101010000110101001110110000101011001000110101000011010100101011000010101") port map( O =>C_1_B_2_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_3_inst : LUT8 generic map(INIT => "0100111101011011101001010010010111110010101100000101101101011010110110101101001001001111010010111010010100100101111100101011000010110000101001000101101011011010000011010100111110100100101001010010010100101101101100001011010001011010110110100000110101001111") port map( O =>C_1_B_3_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_4_inst : LUT8 generic map(INIT => "1001011010010010001101101011011010011011110110011001001010010011100100111001101110010110100100101100100101001001100110111101100100100110001101100110110001101100100101101001011000110110001101101011011010110110001001100010011010010011100100111001011010010110") port map( O =>C_1_B_4_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_5_inst : LUT8 generic map(INIT => "0010010000100000000001000000010000100000001000100010000000100000110111111101111111011011110111111100110101001101110111111101110100000100000001000100110001001100001001000010010000000100000001001111101111111011111110111111101111011111110111111101101111011011") port map( O =>C_1_B_5_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_6_inst : LUT8 generic map(INIT => "0000010000000000000001000000010000000000000000000000000000000000110111111101111111011111110111111100110101001101110111111101110100000100000001000100110001001100000001000000010000000100000001001111111111111111111111111111111111011111110111111101111111011111") port map( O =>C_1_B_6_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 
C_1_B_7_inst : LUT8 generic map(INIT => "0000010000000000000001000000010000000000000000000000000000000000110111111101111111011111110111111100110101001101110111111101110100000100000001000100110001001100000001000000010000000100000001001111111111111111111111111111111111011111110111111101111111011111") port map( O =>C_1_B_7_out, I0 =>  C_8_out, I1 =>  C_9_out, I2 =>  C_10_out, I3 =>  C_11_out, I4 =>  C_12_out, I5 =>  C_13_out, I6 =>  C_14_out, I7 =>  C_15_out); 

C_2_B_0_inst : LUT8 generic map(INIT => "0101100101101001100101101001101010011010011010011000011010011010011010010110010110011010010110010101100101100001100101100001100110011110010110011010011010010110100101100001100101100101100101100001100101101001100101101001101010011010011010011010011010011110") port map( O =>C_2_B_0_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_1_inst : LUT8 generic map(INIT => "0011101111010100101111010100011010111001110101001011110101000110110101000010001101000110001110111100010000100011010000100011101101000010001110110110001010111101010000100011101100100011101111010011101111010100101111010100011010111001110101001001110101000010") port map( O =>C_2_B_1_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_2_inst : LUT8 generic map(INIT => "1010001010011001001001101001101100100010100110010010011010011011011001101011101001100100101000100110011010111010011001001010001010011011010111011011101111011001100110110101110110111010110110011010001010011001001001101001101100100010100110010010011010011011") port map( O =>C_2_B_2_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_3_inst : LUT8 generic map(INIT => "0011110011100001110001110001110011000011000111100011100011100011011110001100001110000111001111001000011100111100011110001100001100011100011000011100001100011110111000111001111000111100111000010011110011100001110001110001110011000011000111100011100011100011") port map( O =>C_2_B_3_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_4_inst : LUT8 generic map(INIT => "1111001111001101110010110010110000110000110100111111001111001111010011000011000000110100111100111100101100001100010011000011000011010011010011011100111100101100001100001101001111110011110011010000110000110010001101001101001111001111001011000000110000110000") port map( O =>C_2_B_4_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_5_inst : LUT8 generic map(INIT => "0011001100000001000000111100000000110011000100110011001100000011100000001100110011001000110011000000001111000000100000001100110011101100011111101111110000111111110011001110110011001100111111100011111100110011001101110001001111111100001111110011111100110011") port map( O =>C_2_B_5_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_6_inst : LUT8 generic map(INIT => "0011001100000001000000110000000000110011000100110011001100000011000000000000000000000000000000000000001100000000000000000000000011111111011111111111111100111111111111111111111111111111111111110011111100110011001101110001001111111111001111110011111100110011") port map( O =>C_2_B_6_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 
C_2_B_7_inst : LUT8 generic map(INIT => "0011001100000001000000110000000000110011000100110011001100000011000000000000000000000000000000000000001100000000000000000000000011111111011111111111111100111111111111111111111111111111111111110011111100110011001101110001001111111111001111110011111100110011") port map( O =>C_2_B_7_out, I0 =>  C_16_out, I1 =>  C_17_out, I2 =>  C_18_out, I3 =>  C_19_out, I4 =>  C_20_out, I5 =>  C_21_out, I6 =>  C_22_out, I7 =>  C_23_out); 

C_3_B_0_inst : LUT8 generic map(INIT => "0101000101011001010110100101101001010101010101010101100001011000101001011010010111100101011001011010011110100111101001011010010110100111101001111010010110100101101010101010101010100101101001010101101001011010100010101000101001011000010110000101101001011010") port map( O =>C_3_B_0_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_1_inst : LUT8 generic map(INIT => "1001011010011110100111001001110001101001011010010110000101100001110001101100011010000110100001100011100100111001001110010011100111000110110001101100011011000110001111000011110000111001001110010110001101100011111000111110001110011110100111101001110010011100") port map( O =>C_3_B_1_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_2_inst : LUT8 generic map(INIT => "1101101111010011110100111101001110110010101100101011001010110010110010111100101111001011110010111111001011110010111100101111001000110100001101000011010000110100000011000000110000001101000011011011000010110000001100000011000000101100001011000010110000101100") port map( O =>C_3_B_2_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_3_inst : LUT8 generic map(INIT => "0100011001000110010001100100011010011001100110011001100110011001101010011010100110101001101010010110011001100110011001100110011010011101100111011001110110011101011010100110101001101011011010110110011001100110011001100110011010010101100101011001010110010101") port map( O =>C_3_B_3_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_4_inst : LUT8 generic map(INIT => "1001010010010100011010110110101100101101001011011101001011010010001111010011110111000010110000100100101101001011101101001011010011010110110101100010100100101001101111001011110001000010010000101011010010110100010010110100101100101001001010011101011011010110") port map( O =>C_3_B_4_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_5_inst : LUT8 generic map(INIT => "0001100000011000011100110111001100110001001100011110001111100011001100010011000111110011111100110111001101110011110001111100011100011000000110000011000100110001001100000011000001110011011100110011100000111000011100110111001100110001001100011110011111100111") port map( O =>C_3_B_5_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_6_inst : LUT8 generic map(INIT => "0001000000010000011100110111001100110001001100011111001111110011001100010011000111110011111100110111001101110011111101111111011100010000000100000011000100110001001100000011000001110011011100110011000000110000011100110111001100110001001100011111011111110111") port map( O =>C_3_B_6_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 
C_3_B_7_inst : LUT8 generic map(INIT => "0001000000010000011100110111001100110001001100011111001111110011001100010011000111110011111100110111001101110011111101111111011100010000000100000011000100110001001100000011000001110011011100110011000000110000011100110111001100110001001100011111011111110111") port map( O =>C_3_B_7_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out, I6 =>  C_30_out, I7 =>  C_31_out); 

C_4_B_0_inst : LUT8 generic map(INIT => "0101101001011010010110100101101010100101101001011010010110100101101001011010010110100101101001010101100011100101010110001110010101011010010110100101101001011010101001011010010110100101101001011010010110100101101001011010010101011000011001010101101001110001") port map( O =>C_4_B_0_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_1_inst : LUT8 generic map(INIT => "0110001101100011100111001001110011000110110001100011100100111001110001101100011000111001001110011001110000111001011000111100011010011100100111000110001101100011001110010011100111000110110001100011100100111001110001101100011001100011010001101001110010111101") port map( O =>C_4_B_1_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_2_inst : LUT8 generic map(INIT => "0001101000011010100001101000011001100001011000010101100001011000011000010110000101011000010110001000011010100111111001010110000101111001011110010001101000011010101001111010011101100001011000011010011110100111011000010110000100011010000111101000011010100111") port map( O =>C_4_B_2_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_3_inst : LUT8 generic map(INIT => "0110110001101100000101110001011101110110011101101001000110010001100010011000100101101110011011101110100011001001011101100111011010010001100100010110110001101100110010011100100101110110011101100011011000110110100010011000100110010011100101111110100011001001") port map( O =>C_4_B_3_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_4_inst : LUT8 generic map(INIT => "1000000010000000000101110001011101110111011101111110111011101110111111101111111010000000100000000000000000000001011101110111011100010001000100010111111101111111111111101111111010001000100010001100100011001000000000010000000100010011000101111111111111111110") port map( O =>C_4_B_4_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_5_inst : LUT8 generic map(INIT => "0000000000000000000101110001011110001000100010000000000000000000111111111111111111111111111111110000000000000001011101110111011100010001000100010111111101111111000000000000000000000000000000001111111111111111111111101111111000010011000101111111111111111111") port map( O =>C_4_B_5_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_6_inst : LUT8 generic map(INIT => "0000000000000000000101110001011100000000000000000000000000000000111111111111111111111111111111110000000000000001011101110111011100010001000100010111111101111111000000000000000000000000000000001111111111111111111111111111111100010011000101111111111111111111") port map( O =>C_4_B_6_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 
C_4_B_7_inst : LUT8 generic map(INIT => "0000000000000000000101110001011100000000000000000000000000000000111111111111111111111111111111110000000000000001011101110111011100010001000100010111111101111111000000000000000000000000000000001111111111111111111111111111111100010011000101111111111111111111") port map( O =>C_4_B_7_out, I0 =>  C_32_out, I1 =>  C_33_out, I2 =>  C_34_out, I3 =>  C_35_out, I4 =>  C_36_out, I5 =>  C_37_out, I6 =>  C_38_out, I7 =>  C_39_out); 

C_5_B_0_inst : LUT8 generic map(INIT => "1011010110100101111101001011010110100101101011011011010110100101101001011010110110110101101001011010110100101111101001011010110110110101101001011101010010110101101001011010110110110101101001011010010110101101101101011010010110101101101011111011010110101101") port map( O =>C_5_B_0_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_1_inst : LUT8 generic map(INIT => "1100100100110110001101111100100111001001001111100011011011001001110010010011111000110110110010011100000100111100001101101100000111001001001101100001011111001001110010010011111000110110110010011100100100111110001101101100100111000001001111000011011011000001") port map( O =>C_5_B_1_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_2_inst : LUT8 generic map(INIT => "0011001011111011111110111100110100110010111100111111101111001101001100101111001111111011110011010011001011110011111110111100110111001101000001000010010000110010110011010000110000000100001100101100110100001100000001000011001011001101000011000000010000110010") port map( O =>C_5_B_2_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_3_inst : LUT8 generic map(INIT => "1010010110100101101001011001011110100101101001011010010110010111101001011010010110100101100101111010010110100101101001011001011110010111010111100101111001011010100101110101011001011110010110101001011101010110010111100101101010010111010101100101111001011010") port map( O =>C_5_B_3_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_4_inst : LUT8 generic map(INIT => "1111010111110101000010100010101011110101111101010000101000101010111101011111010100001010001010101111010111110101000010100010101000101010101010110101010001010000001010101010101101010100010100000010101010101011010101000101000000101010101010110101010001010000") port map( O =>C_5_B_4_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_5_inst : LUT8 generic map(INIT => "0000010100000101000011110000111100000101000001010000111100001111000001010000010100001111000011110000010100000101000011110000111100001111000011110101101101011111000011110000111101011011010111110000111100001111010110110101111100001111000011110101101101011111") port map( O =>C_5_B_5_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_6_inst : LUT8 generic map(INIT => "0000010100000101000011110000111100000101000001010000111100001111000001010000010100001111000011110000010100000101000011110000111100001111000011110101111101011111000011110000111101011111010111110000111100001111010111110101111100001111000011110101111101011111") port map( O =>C_5_B_6_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 
C_5_B_7_inst : LUT8 generic map(INIT => "0000010100000101000011110000111100000101000001010000111100001111000001010000010100001111000011110000010100000101000011110000111100001111000011110101111101011111000011110000111101011111010111110000111100001111010111110101111100001111000011110101111101011111") port map( O =>C_5_B_7_out, I0 =>  C_40_out, I1 =>  C_41_out, I2 =>  C_42_out, I3 =>  C_43_out, I4 =>  C_44_out, I5 =>  C_45_out, I6 =>  C_46_out, I7 =>  C_47_out); 

C_6_B_0_inst : LUT8 generic map(INIT => "0100010001100110001001101011101111011101011001100110011010100010010001000110011000100010101110110101110101100110011001101010101010011001110111010100010001100110100110011101110101010101011001101001100101011101010001000110011010011001110111010100010101100110") port map( O =>C_6_B_0_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_1_inst : LUT8 generic map(INIT => "1011101101000100111110110000000000100010010001001011101100000000010001001011101100000000111111110101110110111011010001001111111100100010110111011011101101000100001000101101110110101010010001001101110110100010010001001011101111011101001000100100010110111011") port map( O =>C_6_B_1_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_2_inst : LUT8 generic map(INIT => "1100110010001000110011001100110000110011011101110011001100110011011101111100110000110011110011001001000100110011100010000011001100110011111011100011001101110111110011000001000111001100100010000001000100110011100010000011001111101110110011000111011011001100") port map( O =>C_6_B_2_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_3_inst : LUT8 generic map(INIT => "1010010101011010010110101010010101101001110100101001011001101001110100101010010101101001010110101011010001101001010110101001011010010110101001010110100111010010101001010100101101011010101001010100101110010110101001010110100101011010101001010010110101011010") port map( O =>C_6_B_3_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_4_inst : LUT8 generic map(INIT => "1010000011111010000001011010000000100100111100100100110100100100000011011010000011011011000001010100111100100100111110100100110110110010010111110010010011110010101000001111101100000101101000000000010010110010010111110010010000000101101000001101111100000101") port map( O =>C_6_B_4_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_5_inst : LUT8 generic map(INIT => "1010000011111010000000001010000011011111000011011111111111011111000000001010000000000100000000001111111111011111111110101111111110110010111111110010000011110010010111110000010011111111010111110000000010110010000000000010000011111111010111111111111111111111") port map( O =>C_6_B_5_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_6_inst : LUT8 generic map(INIT => "1010000011111010000000001010000011111111111111111111111111111111000000001010000000000000000000001111111111111111111110101111111110110010111111110010000011110010111111111111111111111111111111110000000010110010000000000010000011111111111111111111111111111111") port map( O =>C_6_B_6_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 
C_6_B_7_inst : LUT8 generic map(INIT => "1010000011111010000000001010000011111111111111111111111111111111000000001010000000000000000000001111111111111111111110101111111110110010111111110010000011110010111111111111111111111111111111110000000010110010000000000010000011111111111111111111111111111111") port map( O =>C_6_B_7_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out, I6 =>  C_54_out, I7 =>  C_55_out); 

C_7_B_0_inst : LUT8 generic map(INIT => "0110100100011001100101101000011001101001000110011001011010000110011010010011100110010110100101100110100100111001100101101001011011000110011000110110100100111001110001100110001101101001001110011001011011100110011010010111100110010110111001100110100101111001") port map( O =>C_7_B_0_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_1_inst : LUT8 generic map(INIT => "0111000100010001111001111111011110001110111011100001100000001000011100010011000111100111111001111000111011001110000110000001100000001000100011000111000100110001111101110111001110001110110011100001100000001000011100010111000111100111111101111000111010001110") port map( O =>C_7_B_1_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_2_inst : LUT8 generic map(INIT => "0001011110001000100100010110111001100110100110010111011010011001111010000101011101101110100100011001100101100110100010010111011010011001011001101110100001010111100100011110101010011001011001100111011010011001000101111110100001101110100100010110011010011001") port map( O =>C_7_B_2_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_3_inst : LUT8 generic map(INIT => "0110100111100001111010011000011110000111000111101001011100011110100000011001011010000111000101100001111001111000000111100110100011100001100001111000000110010110000101100111110000011110011110001001011100011110100101100111111001111000111010010111100011100001") port map( O =>C_7_B_3_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_4_inst : LUT8 generic map(INIT => "1110011101100111011001110110000110011110100001101000111010000110100110001000111010011110100011100111100100011001011110010001100101100111011000010110011101110001100011101110011010000110111001101000111010000110100011101110011000011001100110000001100110011000") port map( O =>C_7_B_4_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_5_inst : LUT8 generic map(INIT => "0100010101000101010001010100010111011011110110111101101111011011001000100010010000100100001001000101110101011101010111010101110101000101010001010100010101010101110110111011101111011011101110110010010000100100001001000100010001011101110111010101110111011101") port map( O =>C_7_B_5_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_6_inst : LUT8 generic map(INIT => "0100010101000101010001010100010111011111110111111101111111011111000000000000010000000100000001000101110101011101010111010101110101000101010001010100010101010101110111111111111111011111111111110000010000000100000001000100010001011101110111010101110111011101") port map( O =>C_7_B_6_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 
C_7_B_7_inst : LUT8 generic map(INIT => "0100010101000101010001010100010111011111110111111101111111011111000000000000010000000100000001000101110101011101010111010101110101000101010001010100010101010101110111111111111111011111111111110000010000000100000001000100010001011101110111010101110111011101") port map( O =>C_7_B_7_out, I0 =>  C_56_out, I1 =>  C_57_out, I2 =>  C_58_out, I3 =>  C_59_out, I4 =>  C_60_out, I5 =>  C_61_out, I6 =>  C_62_out, I7 =>  C_63_out); 

C_8_B_0_inst : LUT8 generic map(INIT => "1111000000111100111100000011010000001111110011110000110000001111111100000011110011110000001111000000111111000011000011111100111100001111110000110000111111001111111100101011000011110011111100000000111111000011000011111100001111110000001101001111000000110000") port map( O =>C_8_B_0_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_1_inst : LUT8 generic map(INIT => "0011110000000011110000111111110011001100001100110011001111001100001111000000001111000011111111001100110000111111001100111100110011001100001111110011001111001100110000010111110000111111110000111100110000111111001100111100000011000011111111000011110000000011") port map( O =>C_8_B_1_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_2_inst : LUT8 generic map(INIT => "0000110011110000001100001111001111000011000011110000111100111100000011001111000000110000111100111100001100001111000011110011110000111100111100001111000011000011110011110000110000001111001100000011110011110000111100001100111111001111000011000000110011110000") port map( O =>C_8_B_2_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_3_inst : LUT8 generic map(INIT => "1010011001010101010101011010101001100101010110100101101010100110101001100101010101010101101010100110010101011010010110101010011010100110010101010101010110011010011001010101100101011010101010101010011001010101010101011001101001100101010110010101100110101010") port map( O =>C_8_B_3_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_4_inst : LUT8 generic map(INIT => "0110110111000011001111000110100111010011001101101100100110010010100100100011110011000011100101100010110011001001001101100110110101101101110000110011110001001001110100110011010011001001100101101001001000111100110000111011011000101100110010110011010001101001") port map( O =>C_8_B_4_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_5_inst : LUT8 generic map(INIT => "1000010110101001100101011000000110101001011010001010000111101000000101111001010101010110000101111000010110100001100101111000010110000101101010011001010110100001101010010110101010100001111010000001011110010101010101100001011110000101101000011001010110000001") port map( O =>C_8_B_5_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_6_inst : LUT8 generic map(INIT => "0000010100000001000101010000000100000001100000000000000100000000000101110001010101010111000101110000010100000001000101110000010100000101000000010001010100000001000000011000000000000001000000000001011100010101010101110001011100000101000000010001010100000001") port map( O =>C_8_B_6_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 
C_8_B_7_inst : LUT8 generic map(INIT => "0000010100000001000101010000000100000001000000000000000100000000000101110001010101010111000101110000010100000001000101110000010100000101000000010001010100000001000000010000000000000001000000000001011100010101010101110001011100000101000000010001010100000001") port map( O =>C_8_B_7_out, I0 =>  C_64_out, I1 =>  C_65_out, I2 =>  C_66_out, I3 =>  C_67_out, I4 =>  C_68_out, I5 =>  C_69_out, I6 =>  C_70_out, I7 =>  C_71_out); 

C_9_B_0_inst : LUT8 generic map(INIT => "0010000000110011000000000011001100000000001100110000000000110011001100111111111100100000001100110011001111111011000000000011001100000100001000101100110000000000010011000000000011001100000000000000000000110011000001000010000000000000001100110100110000000000") port map( O =>C_9_B_0_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_1_inst : LUT8 generic map(INIT => "0100011001010101100110011010101010011001101010100110011001010101010101011001100110111001101010101010101001100010011001100101010101100110010001001001100110011001100110011001100101100110011001100110011001010101100110011011100110011001101010100110011001100110") port map( O =>C_9_B_1_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_2_inst : LUT8 generic map(INIT => "0010110111000011010010111001011001001011100101101101001000111100110000111011010010010100011010011001011000101001001011011100001100101101110100100100101110110100010010111011010011010010001011011101001000111100101101000110101110110100011010010010110111010010") port map( O =>C_9_B_2_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_3_inst : LUT8 generic map(INIT => "1101111100001100000001001011001000000100101100101111001011001111111100110100111101001111001001000100110100100100001000001111001100100000111100101111101101001111111110110100111100001101001000000000110100110000101100001101101110110000110110111101111100001101") port map( O =>C_9_B_3_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_4_inst : LUT8 generic map(INIT => "1001100110011001100110010010101101100110110101001001010010011001100101011001100110011001101110010110011001000110010001101001010101000110100101001001110110011001011000100110011001100110010001100110011001010110110101101001110100101001011000100110011001100110") port map( O =>C_9_B_4_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_5_inst : LUT8 generic map(INIT => "0001000100010001000100010011001110001000000110000001100000010001000110010001000100010001001100011000100010001000100010000001100101110111111001111110111011101110011100110111011101110111011101110111011101100111111001111110111000110001011100110111011101110111") port map( O =>C_9_B_5_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_6_inst : LUT8 generic map(INIT => "0001000100010001000100010011001100000000000100000001000000010001000100010001000100010001001100010000000000000000000000000001000101110111111101111111111111111111011100110111011101110111011101110111011101110111111101111111111100110001011100110111011101110111") port map( O =>C_9_B_6_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 
C_9_B_7_inst : LUT8 generic map(INIT => "0001000100010001000100010011001100000000000100000001000000010001000100010001000100010001001100010000000000000000000000000001000101110111111101111111111111111111011100110111011101110111011101110111011101110111111101111111111100110001011100110111011101110111") port map( O =>C_9_B_7_out, I0 =>  C_72_out, I1 =>  C_73_out, I2 =>  C_74_out, I3 =>  C_75_out, I4 =>  C_76_out, I5 =>  C_77_out, I6 =>  C_78_out, I7 =>  C_79_out); 


out_fin <= C_0_B_7_out  & C_0_B_6_out  & C_0_B_5_out  & C_0_B_4_out  & C_0_B_3_out  & C_0_B_2_out  & C_0_B_1_out  & C_0_B_0_out  & C_1_B_7_out  & C_1_B_6_out  & C_1_B_5_out  & C_1_B_4_out  & C_1_B_3_out  & C_1_B_2_out  & C_1_B_1_out  & C_1_B_0_out  & C_2_B_7_out  & C_2_B_6_out  & C_2_B_5_out  & C_2_B_4_out  & C_2_B_3_out  & C_2_B_2_out  & C_2_B_1_out  & C_2_B_0_out  & C_3_B_7_out  & C_3_B_6_out  & C_3_B_5_out  & C_3_B_4_out  & C_3_B_3_out  & C_3_B_2_out  & C_3_B_1_out  & C_3_B_0_out  & C_4_B_7_out  & C_4_B_6_out  & C_4_B_5_out  & C_4_B_4_out  & C_4_B_3_out  & C_4_B_2_out  & C_4_B_1_out  & C_4_B_0_out  & C_5_B_7_out  & C_5_B_6_out  & C_5_B_5_out  & C_5_B_4_out  & C_5_B_3_out  & C_5_B_2_out  & C_5_B_1_out  & C_5_B_0_out  & C_6_B_7_out  & C_6_B_6_out  & C_6_B_5_out  & C_6_B_4_out  & C_6_B_3_out  & C_6_B_2_out  & C_6_B_1_out  & C_6_B_0_out  & C_7_B_7_out  & C_7_B_6_out  & C_7_B_5_out  & C_7_B_4_out  & C_7_B_3_out  & C_7_B_2_out  & C_7_B_1_out  & C_7_B_0_out  & C_8_B_7_out  & C_8_B_6_out  & C_8_B_5_out  & C_8_B_4_out  & C_8_B_3_out  & C_8_B_2_out  & C_8_B_1_out  & C_8_B_0_out  & C_9_B_7_out  & C_9_B_6_out  & C_9_B_5_out  & C_9_B_4_out  & C_9_B_3_out  & C_9_B_2_out  & C_9_B_1_out  & C_9_B_0_out ; 
cor_out <= cor_in;
end Behavioral;

