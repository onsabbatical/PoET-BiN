--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   01:13:09 07/28/2019
-- Design Name:   
-- Module Name:   D:/siva/Masters/Thesis/07_ETE_19/part_svhn/mnist_tb.vhd
-- Project Name:  part_svhn
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: minst_check
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY mnist_tb IS
END mnist_tb;
 
ARCHITECTURE behavior OF mnist_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT minst_check
    PORT(
         inp_feat : IN  std_logic_vector(511 downto 0);
         out_fin : OUT  std_logic_vector(79 downto 0);
         cor_in : IN  std_logic_vector(79 downto 0);
         cor_out : OUT  std_logic_vector(79 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal inp_feat : std_logic_vector(511 downto 0) := (others => '0');
   signal cor_in : std_logic_vector(79 downto 0) := (others => '0');

 	--Outputs
   signal out_fin : std_logic_vector(79 downto 0);
   signal cor_out : std_logic_vector(79 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: minst_check PORT MAP (
          inp_feat => inp_feat,
          out_fin => out_fin,
          cor_in => cor_in,
          cor_out => cor_out
        );

   -- Clock process definitions
   --<clock>_process :process
   --begin
		--<clock> <= '0';
		--wait for <clock>_period/2;
		--<clock> <= '1';
		--wait for <clock>_period/2;
   --end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

     -- wait for <clock>_period*10;
inp_feat <= "00000000000111111011111011111111111111101110110000000111111111101111011101111001011011011111111100000000011111111111111111111011011001001111111101100111111111110111111111111111111111101110110000000000011111111111111100110011111011001000000111101111000110111111111111111110111111101111100011111010100011111110110001111111001011101111010011101110111001110010010111110011111111111000111100110111100011111111111111111101100111111111011111110111010111111110111011110111111111101111000011111111111101111111111001011111";cor_in <= "10011110101010111001100110100100101101011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11111100000001100001000000111110011111111111011111101110000101110000111110111011111100100111011111110000000000011011111111111111111100010000010111110111101111101001101011111111000000010111111011111110000000111111111111101001011101111110110111111111110110011110111111111011000000111111111111110111110111011111111011111011000100010011011111111111111111110111000010100111111111111111110011111111111111011101111111111101111111011111111111111110111100111111011101010111011111111111001111110001111110111111111111110111";cor_in <= "10011110101010110100010010011110101101011000000010111000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00000000000000000111011111111110111110111110011000000000000000001010101111110111001001100000110000000000000000000001011111101110001100100010011001111010111011001110111111111111000011111110111001100000000000001111111111011011001111101100110011111110111011100111000100010011011110111110111011101111110011001110110011101000111101101110111010111110110011100011001001100100111111111111011111110100011001101111111111111111111110110011001111101011001100110110011011101110011101101110111011111111111110110110111011101100";cor_in <= "11110111010001101001100110011110101111001000000010101011101000001001011110000001" ; wait for 10 ns; 
inp_feat <= "11111100010001100011101111111111001111111101001100101110110011001101111101111111011111001111111001110000110111100011110111110111011111001100011111111111110111101100111010001111111011001111011101110011111011101111011101111001111110110111111111111111111110111100111010000001110011011111011110111111111011111111011001101111001111111111011101111111001100111111110111000010111110111101011101111110100111111001011101111001111111001100000011110100010011111111001111101111111100110111010111111100011101111111111111010010";cor_in <= "01001100101010111001100110011110101101011001011110100101101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "01110111000000001111110011101111111111101111110101110110011101010011011111111111011111111000101111110111000010000111101111111111011101110101111111101111101101011011110011001111101001101001111111111111101100001011111111110111010011111011001010011111111111111111110011100111111001001111111111001111111111111111111111111010111111001101111111111111111111111111001111001000110011111111111111101111111111111111110111011111111100111100000011111111010000011111111111110111111011111111010111111111111001111111111111011101";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "01000000000000000111111110111111101111111110011000000000000000001001100110110011001001100100110000000000000000000101111111101110001100000000010001100010010000001111111111111111000011111110111001100000000000001111111111111011011101101100110011111110111001100101000100011111001110111111111011101111111011001110110011001000001110100110011011111110010001000111000001100100011101111111111110111000001011101111111111111111101110110011001111001001100100110110011011101110011001101100100011111111111111110111111011100110";cor_in <= "11010001010001101001100110011110110000111000100010101011101010101000110110000001" ; wait for 10 ns; 
inp_feat <= "11000011111100001011111111101111111001101110111111110111011101111111111101111111111101111111101101000111011100001111111111011111011001111111110111110111111111111101111111011111101011101110111101111011011101111111100110011111011011001111101111111001110111111001111011101111111111111100111111001100111111111110111111110000001111110100110101111111111111110111111100110000111111001001111111111000011111111111111111011101111111110010000011011111111100000110111111111011111111111011111111111111111111001100001111111101";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110111011001111101111111111111010001110011000111111101111111101111110011011111011101110100011011111111111111101110011101011111111101110111001101110111111001111011000011001111000001101111101111011111111111100011001110011101000011111111011101011011101111000011001011001101111011101111101111001111111111111011001000111110111111110111000101111011000100111111111101110000111111110101001111101011111111111111101110011100111111001000000111110111000011000111111101110111111011111111000101110111100000011111111101100000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110100000111" ; wait for 10 ns; 
inp_feat <= "11111111001011111111111100000011001101100100000111111110111111100001111111110001011111011111111111111111110111110011110111111111111111110011111111111111111111011001111011111011111010100001001111111111111111100011100111111111001000010011111100111101111101111001110011101111111110000001110110000111001100110111111111111111011100001100110000110111111110111111001111001110111100010011000101111111111101110011110011111111111110011110111011111111110011111111011100111110001100111111110011111011110011101101001100101101";cor_in <= "10011110101010111001110110011110101101010010011010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00000011111111110011111111101110001101111100111100110011111011101011110101111111011111111111111000110011111111111111111111011111001001111111111111111110111111111111110111001111011111101100111100010011111111001111100100110011111011011111011011111001000111111101111111101111111111111101000011001000011100111100101101111111011101111111000011111011001101111111111111111000111111101101010110110111111111111111111100110111111111111110011111001111011111111100101111111100111010110111000111111111111100001101111100000000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 
inp_feat <= "11110000100011000011111010111111111111111101010111101110110111101111111111111001111010001111111101110001100011101101111111011111111110001001111111111011001111001100111011111011110010001001111101110011001011111111011101110111110110110011011111111111111100111111111000000000100010011101111111111011101101111111001000101111000011011111111111111111111100111111110011011110101111111111100101111111110111111111111111110111011111001101110011110110000011001111101110111110101101110111011111110111111111111111111110110001";cor_in <= "01001100101010111001111110011100101111001000000010101011101010101000110110000001" ; wait for 10 ns; 
inp_feat <= "11111110111011000011111110111011001111111111011101111110101111011101111111111101111110001110100001110111110011001111101111111111111111111111110111111111001101111110100011011111111011001111111101110111111010011111001101100111111111110111101101111111011111111100110011001110110111111111011111111111011101110111011011101111011111111111001111111111011111111111111110000001111110111011011111111111111111110011111011001111111110001000110111111110110011001111111111110011101111110111001111110100111100011111110100011011";cor_in <= "10011110101010111001100110011110101101011000000001000000101111101000110110000001" ; wait for 10 ns; 
inp_feat <= "00110111011011111011111111001110011101110101111101110101111011001111010001111111011111111110111001110011011111101110111111111111001101111111111101100111111111101011110011001111111011101101111100110011011101101101101111010011110011011111011011011011011000110011111011001111111011101111111111001111011100111011111111111111011101111111000011111111111111110111111111101000010111111111010111100111111111111111111110110001111111001100111100101111001011111111111111110110111011110111001111111111001001011111111101000000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 
inp_feat <= "11110000010001101111110111111111111111001101001101111110110011001111011101111101110111001110011101110001110011101111110110010111111110001100111011110001110111001100101001111111100011001111011101110011011011101111011101110011101100110011011011111111111110111100100000000001110111011111111111111111111111110111001000000110111111011111111111111110110100111111110111101100111111111111110101110110110011101101111101110111100110001000000111110100000000010111101111101110101101111111100111011110111111111111111111010001";cor_in <= "01001100101010111001100110011110110000001011000010101011110001001000110110000001" ; wait for 10 ns; 
inp_feat <= "01100000000000001111111111111111011101100110011000100010001010101000101010101011011000000100011001100101000101010011011001010111011100000000001011110010001000001011111111111101110011001100110001100100000001101111111111011011001001100100001011111110111011101111000100010001011101110111111111101110111011100110111011101010111011101110111011111100110000000111011001100110111111111111111110111011100011111110111111111111111101110011001111110010001000110110001001100110010001100110011011111101101110111110111001100110";cor_in <= "10011110010001101001100110011110101101011000000010101011101000001000110110101001" ; wait for 10 ns; 
inp_feat <= "11111110111111011111110011010011111011110001001111111111111111111111111111011111110111110111111111111111111111111101111011111111111111001111011111111111111111101111111111100110100010000000000011111111111111110111011101111111100100010111111111111111101111111111111111001111100011101001110101110000000100000111111111111111110011110011011111111111011111111101111101111111111111100011101111111111110111111111111100011111111111110111111111111111111111111100111111111111001101110011111100000111011111111000111100110011";cor_in <= "10011110101010111001100110011110101101010011110010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00110111000001111111101111111111011101101110110101110111011111101011011011110111011111111100111100110111101111110111111110011111001101111101011111100111111011101111110011101111111011101101111110110011011111111011101111110011110011011011001111011111011110110111110011101101111111001111111111001111111101111111101110110111011101011111110111111111111101111111101111111110111111111111010111000011111111101111110111111110111110111101110001111111000011101111111111110110111011110111001111111111001001111011111111000000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 
inp_feat <= "00000000010111110011111011111111011111101100100000000111111111100101111101111100011011101111111100000000111111111111111011101011011001001111111111101111111111111111111111111111111011101100000000000000011111111111100100000011110011000000000011101111000010001111111111101111111111001111000010101010000001101111110001111111011011101111000011101110111001111010111111110011111111111100101100010111100011111111111101111101101111111111011111110111111111111100100011110111110010100011000011111111111101111110111011011101";cor_in <= "10011110101010111001100110100100101101011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111111100111111111110111111110111110011000011111111111111111111111111001111111111111111001111111111111101111011111101111111111111111111011111111111111111101110101110101110100010000010000111111111111111110111011111111100000101111111111111011111101111111100111111011100110000010010100101100001011100111111111111011011111110110011000111100111011111001111111101110010111111000111001111111111111111111111111110011000111011111111110011111100111011101111111111110011010101111001000111110111001100001001111101110000";cor_in <= "10011110101010111001100110100100101101011110010010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00101111111100001110111011111111011011101101011111110111111101000111110011111111111101111100001011111111011001010010111111111111010101110111000111111111011100001101110111001011011011101001111011011111111100001111101111111100010011011111100011011011111111110011111111110011011011100101111111001111111111000111111111111111111101101101111101111111111111111111111100011000111111011111111111110001111111111111001111011111111111111111100110111111010000111101111111111100111111111111000111111111000001011101111111000100";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001001011110000001" ; wait for 10 ns; 
inp_feat <= "00100011011111100111001011011110101101110111001100110111010010001111011101111111011101111111111000000011011111101111111100010111001000111111111001110110111111111111111101001111011011101111111100110011011101001111100110110001111011111111011011111001000101001111111111111111111111101111111011101100101100111110111100111111001101111111000011101111001101111011111111011000011111001111011111110101001111111111111110010001111111111001001110001111111111111110111111110100111111111111001111111111111100011110101110100000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 
inp_feat <= "11110111111000000111111111010101010101110011011111111110111101000101111111111111111111101100011001111111111101001011011111111111111111110111001111111100011101101100110011011110110011000000001101110111111010001111001110111111111100110111011101111111111111111100110011100100110110110001011111100110011101110110011011101110111111110001011111110000011111111111111100001100111111011011111101111111110110010011000111111111111011001100110011111100110111001111111101110111101001110111111111110101000111111111001101110111";cor_in <= "10011110101010111001100110011110101101011110001101000000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111110011000011111111111111001111111110011100111110101011011011111111111101111110011100100111110011100111000111111111111111011111111100110111101111001100111001100011001111110011001110111111110111011110001111111101110110111011111111101101111111111111111010110000001110111011011111111111011111111101111111001111001110011111111111001111111111011001111111101110010001111111111001011100111111111111111111000100011101111110010000100011100110100011001111111111110011111001110111001111111001011000111111111100110101";cor_in <= "10011110101010111001100110011110101101011000000000011001101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "11111111111011101111111001011111011111110011001101111111111111000111110011110101111101111100111011111111111011111110111110011111111111110111101011111111111110001111110011001111111011100001011100110111111011111111001111111111110000110111111000111011111101111111111110011000111011000011111110110110011000110111111111111110011000001111111111110111111111111111011110111100111101111111000111111111111111100111101111111111111111111111110111111111100011001101011100111111100000110111111111110011000111110111011101110011";cor_in <= "10011110101010111001100110011110101101010011110010101011101111101000110110000001" ; wait for 10 ns; 
inp_feat <= "00111111011000001110111011111111011011101111001111111111111101000111010011110111111111110101101111111111010001000110111101110111010101110101010111111111001101000011100010011111011011101000011111110111111100011001101111111101110000110111000010111111111111110011111010110010111011000111111111001111111111101111111100011111111111001111111111111111111100111111011101010100110111111111011011111111111111111111010111011011111100110111000010011111000000011111111111110011111111111111001111110111001001111011111111010001";cor_in <= "10011110101010111001100110011110010110011000000010101011101001111000110110000001" ; wait for 10 ns; 
inp_feat <= "11111110000011110001110111111111000111111101101100101110111011100110111111111011111011001001101101110111110111111001110011101111111111011011111111111111111110010000111011101011111011101111111111110001011011101011011101100111111111110011011101111110111101101100111011100001110110011101111010111111111101011111101001111101111110011111110111111111111101111111100111101110111110111110110101111110110101111100011011100101111111101110100111111110110011011111101111111101111110110011000111111110111011001011111111011100";cor_in <= "01001100101010111010001110011110101111001000000010100101101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00000001011111111110110011001111111011001100000101000111011111110111011100001110110011111111111100000001111111111110111011111111010000001101011111001111101111111111111110011111111011001111001000000000111111111001100100111011110010000011001011001100100010110011001010110111111011101111111011001100100000111100100101111111111011111111110011001111001100111100111111110001111111101100101101110111111011111111111101111111111111111111111100110001001111111100110001110100111011111111000011110111011101111100110011010000";cor_in <= "10011110101010111001110010100100101101011000000010101011010001011000110110110101" ; wait for 10 ns; 
inp_feat <= "10111111011100001111111011001111111011101101011101110111011101010111000011111110111101110101101001110111001010000110101111111111010001110101101111110111001100111111110111011111011011101001111111110111011100001011101111111100010011011111011010011101111011111111111011110111011111000111111111001011111111111111111111110000111111001101111111101111111111111111111111001010111111111111111111110101111110111111000111111001111111110001001100011111001100011110111111111101110011111111010111111111000011011111111111101111";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110000000001111111111111111111111111101111001111100110010111111101111101111110110001001111011101111001110011111001110111110111111100011111111011110011101111101100110100111111110010001111111101110110011011111111111101110001101110110111011011111111111110111100110000010011100011011111111111111111110010010111011001101101110111111111111111111111001100011111110111101111111111111111111011111111001010111101111111110001111111011100110011100100000010111111011101111111001111111011100111010110111101111111111111010011";cor_in <= "01001100101010111001110011000111101101011000100010101011101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "01100000001000111110111111101111101001100111011110100010101100111011101010111010001000100110011001100101011111110010011101110111011000000011001011100100011101001001111111001101000001100100011001100001010000011111100111011101001001000100010011111111111111111001000100011001011001110111111111001110111011100110101010001101111011111111111100111000101100000111011001100111111111111111111110111101111101111111111111111111011101110111111111110011110010010110001000100011011001110111011111111011101111111110011001100011";cor_in <= "10011110010001101001100110011110101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110110111101110111111100011111011111101011001101110111111101100111001011111110111111111111001100111111111111111110111110111101011111110011011111111100111111110111111110111110111011000010111000110111111100111011001110111001110000101110110000110011110110111111111111011111111011000011111110111100111010010111011111111011011011100111101111110111001110011111111111110111111111110110011001111111101101111111101110111001111111111111111111111110111101111100011001110011100001111111000111101111000100111110111111010111";cor_in <= "10011110101010111001100101011010101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00000000001000001110111111111111001001100110001000100010001011101010101010101010101010100100001011001110011111110010011001100111011000000010001111100100010001001001100111011110000001100110000011000100000001011111100111011101010000000000000011101111111111110011000100010001011001100111111111001100111011101100100010001000111011101111111101000000100000000110011101110110111101111111111111111111111111111111111111111011011101010111101100110011101110010110001000100010111011101110011110111111101110111110011001100110";cor_in <= "10011110010001101001100110011110101101011001011110101011101000001000110110101001" ; wait for 10 ns; 
inp_feat <= "11110110111100111111111000011110011111110001001111111111111101111111010011111100111101110111011111111111111111111111011111111111111101110011011111111110111101101111100110111111110010000010111001111111111100110001001111111001100000111111110101111001110111011111101111111111111010100111111100100100111100010111011111110011111111100011101011110011101110011111111100110111111101101111111011111101111111000111101110011001111111110111111111111111111101110100011101110011001101111111001100010111000100111101111100100011";cor_in <= "10011110101010111001100101011010101111001000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111000000001100110010111111100011011111101111111110110100010000111111111100111111100001101111111111000000100111111011111111111111111001101111111111101101001011110011110111000000000111111111111111000000001111111111101100100110111111000000011111111111111111111101110111101010001111111110011111011011101111111111100110011110001101111111111111111110111111100110010011100110111111111101001111100101111111111111011111111110011111101111111111110100011111111110111001111101111111100111110011110011011011100111111011";cor_in <= "10011110101010111011001011000001010010101000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00110000001011110101011111111111001101110110110000000000011101111111011111111000011001101111111100000000011111111111111111101111001100101111111111111110111111111111111111111111011111111110111000010000011111111111111110010011111011001100100111111011100101110101111111111110111111101111111011011111100000011110111111110111001101101111110010000111011101111111100011111111011111111011100010110111010010111111111111110001101111111111101111111111110111111100110001111111111011001010001011111111111111111111111110111111";cor_in <= "10011110101010111001100111000001101110101000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11111110100011110101000111001100000001111111110011111111111111100010111111110001111111101111111111110000000011110110111111101111111101101101111111111111111111111111111111111011101101111100111111111100000011110111111000010011011111101001011101111111110100011111111111111111000011001111111111011011111010011111111100110111000100001111111111111111111111111111100011111111011110011111100011111111111111110100111111110111110110111111111111111111011101111111110011111111110011110111011111110000111111111001111111011001";cor_in <= "10011110101010110100010010011110101101011000000010101011101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "11001100010011111010100011101111011011110110110010001000011111101010111101111100111011011111111110111100111111111111111111011111111101101111011111111111111111111110111111111111111011101111110111101010011111111111101010010011111011001101001001111110110010111001111111111111111111111111111011111111100000011110111110111111011000001111110011111111111101111110100111110101011101111110010110111111111010111111111110110000101110111111011111111011010111111110111011110111111111110111000011110011011101111110111001010100";cor_in <= "10011110101010110000101010011110101101011000000010101011001110011000110110100101" ; wait for 10 ns; 
inp_feat <= "01000000000000001111111111111111011001100110011100000010001010101010101010101010011001000110001001000101011101110011011001100011011000000000001111000010000001001001101111011111000001000110010001000000000000001111110110111101011001000100000011101110111111111011000100010001011101110111111111001110111011101110101010101000111011101110111111001100000000000111011001100110111111111111111110111001110111111111111111111011011101110111101100110010101110010110001000100010011001100110010011111011101110111110011001100110";cor_in <= "10011110010001101001100111010001101101011000000010101011101000001000110111001010" ; wait for 10 ns; 
inp_feat <= "11111110100000110001111001111110001111111111001011001110001101101111111110111011111010000111011111111000000101011111111111101111111111110001010111111111101111111000111111111100111111111110111101111110000100111111110011011001111101101111111101111110111110011111111111111111110111111111111101111111110011011111111011110011100100110111111111111111111111111011000001110110001111111111111011111111011101111101111111111011100110101111111111101110101100111111011101110111111101111111011111111001101111110110111111110001";cor_in <= "10100110101010110011111010011110101101011000000010101011101000001010011110000001" ; wait for 10 ns; 
inp_feat <= "01100000000000001111111111111111001101110110011000000000000000001010101110110011001000000000010001100010000000000011100111011110001100000000000001100010011000001100110011111111000000001111111001100000000000001111110111011111001001101100110011111110111010101001000110011001001100110111111111101110111011001110110011000100111011111111011000111000100000000111011001100110111111110111011111111101100011101110111111111011111100110111111111111101110000110110011010001010011001100100011011111101110111110110011011100110";cor_in <= "10011110010001101001100110011110101101011011010010101110101000001000110111000101" ; wait for 10 ns; 
inp_feat <= "00000000000000001110111111111111111101100110011000100010001000101111101111111010001000100000000011101010101001100011011101100110001100000010001001100010000000001101110111111101000001100110011001000000000000001111110111011101001000000000000011101110111011100101000100010001001101110111111111101100110011001110110011001000111011101110111011111110111010100110011001100111111111111111111111110110111111111111111111111111111111111111111111111001100110010110011001100110011001100110011011111111101100111110011001100110";cor_in <= "10011110010001101001100110011110101101011000011010101011101000001010011110000001" ; wait for 10 ns; 
inp_feat <= "11001110000011111111111111101110011101101110000111101111011111110010111111110110111011011111111111001111111111111111111011111111111001100101011111001111011011111111111110111111111010001110111011101100011101111111101110011011010011101111000001101111110110111011101110111111111100111111111010001110110010111100111000111111111101111111100011100111111100111110011111111101111111111100011111111111111011111111111111110011101110111111001111111111011111111110111001110111110111110111000011110011011111111110111011110010";cor_in <= "10011110101010111001100111001010101101011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "00110011011000001011111110011111001101110111011100110001011001101111001001111111011101110100111101110011001100010111001110111101001100110111110101110111011000101011110011001111001011101110111111010011001100001101101111111110110011011111000111011011111111110011101010101010011111101111111111001111111111111011101110000010111101100111011111110111011001010111111111011100010111111111111111111001001111111111101111001100111111101100100010101111110000001011111110111111111011111111001111111111110000111111111111111101";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "00111111110001100000101100011110000011111111011011101101111001101110001111110000111111110110010011111111000011000111111111111111110111110110010011111111111010001111101111111111000000110110111011111101110000100111111111101011011111111110100001100111111111101111111111111111011100001110111000011111111111001111111111000000111100010010111011111111111001001111100100101110001001111111111110011111111111111111101111111111111110011101110111111111110100111111111101100110111101101111001011111111001101110111010011111110";cor_in <= "10011110101010110100010010011110101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110110111000010011111010111110011101101111011101100111111100110111100011111011111011101010011100111111111001111111011111111111011111010011011111110100011101100111111111011101111011100000011000110111111000111111101111111101110000100111010000111111111111011111111110010111111011000011111111100010111010100111011111101011011111100111111111110001101111111111111100110111111111111111111001111111111111111011101111111111111111110111111111101111111110111110011001100011111100110111011111111111000100111110011001100011";cor_in <= "10011110101010111001100100101110101110001011000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11100100111011001111111011111111011111110011001101110111111111000111101011101011011111111110111000111111111011101111111111111111111111010111111011111101111111001111111111101111110011000010001100110111111111111111101100111101111100110110010011111111111111111110111100111101111011101111001111110111111100100111011111001110111111111111011111111111001111101111111000111100111111100111101101111111111101111111111111111111111111111011110111100111110111011111011101111111011101110111011111000111111111011100111101100111";cor_in <= "10011110101010111001100110011110101101010011110010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11100010001100111110111111111111011001100111000100101010101111011110111010101111010000000000000011111111011111110110001011111001011001100010001111100100010001001001100111001100000000000100000011001000001101110111111110011101011011000100010111111011101111111011100110011001011001110111011111001100111011100100000010001010111001100111111101100000000000001111011101110011111101110111111111111011110111111011101110111111111111110111101111010011001010110100001000100011110011000110011111111011101110111110111001110111";cor_in <= "10011110010001101001110110011110101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111011101101011011111101110001101110111111011111110011101111000111111110111111101111100111111111111101011111111111111111110111101110111010111111110111101111000011011111011011011111110110011111111011100111111101111001001111111111100000000011111111011111110111011110011111011111110111010111111111111001111111101111001001100011100111111111111110111111111011011001111010111001111111111011111111111110111100011111111111111011111111111111110001100111111111101000110011111010011001111110001000111111011110011111111";cor_in <= "10011110101010110100010010011110101110001000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11000011011100001111110000011111011001101101111101110111011001001111100011111111011101111100100101110111011011100110011110010111000000110111110101111111111111111111100011001111111011101111111101110011011101001111101110110111100010111111011111011001111111101111011111001111111101101101111011001011111101110011011100111000011101101101110101111011011101111111111110111000111111111111101101110001011111111011111100000000111111111111100111111111111110011110111100110111111111101011000111111111111000001101111111111101";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001010100011000011" ; wait for 10 ns; 
inp_feat <= "00111111111000001111110111111111011101011111111101110111011101010111110111111111011111111000000111111111011011010111101111111111011101111110010011101111111100100011110011001011000011101100010110111111011110001011101111111110110011111111000010111111111111110111010011100000111011001101011111001011111110110111111110100001111111001101111111111011111000111111111111011101111111111111110111000011111111111111100101110101111100111001000001111111010000001111111101010111111011110011011111111111000001111011111111111101";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110100100000001111110110010010011111111111011101110111110000000101111111111111111111001110011001111110110000001011111111111111111111010011011011110011001011100100110011110111110011010011111101110110110000001111011111011111111100111110111001111111111111101100110011111111110010110011111111100111111111110111011011101101111011110011111011111111111111101111110000001000111111110111111101111111111001110101100111111111111110011000100111111100110011011111011101111110101101111111111111111101101111111111010111000110";cor_in <= "10011110101010111001100110011110101101011001101101000000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111100111101111111110000111111111011110011011111111111111111111111011111111110111111111111001111111111111111111001111101111001111111110111011111111111111111111111110110011110100010000110111011111111111110111111011100111001100001111110110111111111101110011101111110111111110010000111110011100000111100001111111111110111111110100111000011110110011110111111111101110111111011001111011111111111111110011111111110111001111111111111111111111111111111111111111111010111001101111111000111111111011100111010111110000111";cor_in <= "10011110101010111001100101011010101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110111111111101110111000010111011111110011001101111111111011000111110011110110111101111111111011111111111011101110111111111111111111110111111111111111111111111111110011101111111011000011111101111111111111001011001111111110110100111111111000111011111001111111111111111111111011000011111010110011011101110011011111111111111001111111000001110111111111111111111110011000111100010011000111111111111101110111011111111111111111011100110111111111111011111111011111111100001100111111100111110111110011011111111100000001";cor_in <= "10011110101010111001100110011110101101010010011010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110111111111001111110011010001111011000001001111111111111111101111111111101111110111111111111101111111111111111111111111111111111111110111001111110111111111101011111111000111110011100000000011111111111111110101001100111111100100110111111111101011101111111111111101101110111011101101111111100001001100010111111111110111110111110011010111110111011111111110111100111100111111000011110111111100111111111111111111111111111111111101111011101111111011101110111111111110001101110011111110001111111101111000101100110110";cor_in <= "10011110101010111001100110011110101101010011110010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111110011001111111110100000011110110111111111111110110011101000111111101100111110001100000111111111110010001011101011111111111111111100110111101011101111111110000011111101110010000110001111111111111110001111011111111111101111111111101101111111111111011110100010001110110010110111001111011111011111111111011011101111011111110111000111111110111111111111111110000000111101010001111111111111111011000011011000011111111110000000110011111110110011011111110111110011000011110111011111111000111100111111111100011101";cor_in <= "10011110101010111001100110011110101101011001100101000000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11110000000001101111111111111111111111111111001101100100110111001111111101011111110011111110111001101000100011101001111111110111111110001000111011110011111010001100111110101111110011011111111101100000010011101111111111110011101100110010011011111111111110111100100000000001101111111111111111111110111011101110011101010100111111111111111111111110100000101111111111111110111111111111101111111111110111101101111111110011101110011001100111110000000100011111011101010100101111110110001111010111111101111111111111110011";cor_in <= "01001100101010111001100110011110101101011000000010101011110001001001011110000001" ; wait for 10 ns; 
inp_feat <= "10010111011100001111110101011111011011011111111101110100011000010111010011111101111101110100100111110111011000010110111111101111010101110111100001111111111100111011110011101111011011101000111110110111011100001111101111111110110010011011001011011111111111111011111011110110011111001001111111001011111111110111111101110000111101001101111111111011111111111111111110011001111111111011111111110101111110111111011111111101111111111101101010111111000000000111111100011011111111011011001111111111100011001101111111111111";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001010100010000001" ; wait for 10 ns; 
inp_feat <= "01000000000000000111111111111111001101101110011000000000001000101011101111110011001001100110010000100000000010100111011111101110001100100010010001100010111010001011111111111101000011011110111001100100010000101111111111111001011001101100100011101110111011100101000100110001001111111111111011101100110011001110111011101000111101101110111011101111111011000110011001100110111111111111111111110110011011101011111111111111111111111111111110101000100100110110011011101110111011111110011011111111111101110110111011101110";cor_in <= "10011110010001101001100110011110101101011000000010101011101000001001011110000001" ; wait for 10 ns; 
inp_feat <= "00010111111011111111110111001110111011101110101101110101111111100111010011111111111111111111111001110011111111111110111111111111001100111111011101111111111111111111110011001111111011101101011100010011011111001001101100110010110011010111001011010011011010111111111011101111111111101111000111001011011100111011111101111111111111111111000011111111001100111111111111100100110111111101111101100101111111111111111101110111111111011110011111111111011111111110111101110101111011110111000111111111010000011101111111000000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 
inp_feat <= "00110111011111110111111100001000011100100001011100111111111111101011111111111111011111111111111000101111111111100111110101111111001100110111111101111111110011111111111111011111011100100000110000110011011111101100110101111111000000011111101011111111011111111111101011011111111111101101100001100000000001110011111111111111111111111111000001101101111111110111111111000100111110110000011101111111111111111111111111111111111111111100111110011110111011110011001111101100000101111111001110111101111110010111001100000000";cor_in <= "10011110101010111001100110011110101101010011110010101011101000001000110110010001" ; wait for 10 ns; 
inp_feat <= "00000100011011111110111011100011111011101000000001000111111111110111011101011110110011110111001100001111111111111110110001111101000011001111011111001111111111111111111111111111111011001100000000000011111111111011101100111011100010000000100011001111100011011111011100111111111011100111000011001000000000111000000001111111110011111111000011001000000100111100111111110001111111111100111101100111100011111111111101111110111111111111111100110101111111110000010001110111100010100001000010110111011100111110110010000001";cor_in <= "10011110101010111010100110011110101101011001100110101011010001011000110110110000" ; wait for 10 ns; 
inp_feat <= "01110111110111101000101111111100001001111111110001111111111111101000111111111111011111111100111000110111111111110101111111011111011101111111111111111111111011111000111111111101010001111110101101110111011111101111110111010111011111111111011110010011011101101110111111011101111011111101101111011001011001110011110110111111011111101111101111111111111101111111111011111100010101111011000010111111111111101111110110111100111111101001100011111011111111001111111110111111111111010111011111111100100011111110011111111000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000000011111110000001" ; wait for 10 ns; 
inp_feat <= "00110011000001101111111111111111011101111111000001110111111111101111011111111001011101111100111011110111111111110111011111011111001101110101011101100111111011101111110011101110011001001000000110110011011001111011111111001111000001110001000110011111111101110111000011001100011011111111100111101111111001101011101011111111111101111111011111110111010111111111011110111100111101110111100011111111111100101111100111111111111100111101110000110111110111101111101100111111111101111111001111110111011111111111011100111100";cor_in <= "10011110101010111001100110011110101101011010110110101011101000001000110111011101" ; wait for 10 ns; 
inp_feat <= "01110011111101101011111111111110101001111110011101111111111111111111011001111111011101111111011001110111111111111101101111011111011101101111111011111110111111001111010111111111111011101100110000110011011111111111101110011011111111011101000011111111011111111111111111111011111011101100101011111100111100000011111110110111011111101110111011111111011100001111111111101110110101001111011111111011011111111101111111111111111111101111111111111111111111111111111111100110110111010111000111111110011100111110111111001111";cor_in <= "10011110101010111011111001011010101101011000000010101011110001001010011110000111" ; wait for 10 ns; 
inp_feat <= "00101111111111110111111111011111001101111111111111111111111111111111010111111000111111111111111111011111111111110111111111011111101111111111111111111110111111111111011111111111011101111100100011001111111111111111110100010011011011001100000011110011011011101111101111111111111101101101100000001000111111101101111101111111111101111111000011111101111111111111111111111101110110101011111110100111110111111111110111110000111111011111011110111111111011111100111111111111110111011011001111111111011101111001101101011111";cor_in <= "10011110101010111001100110111110101101011000000010101011010001011000110110100101" ; wait for 10 ns; 
inp_feat <= "00100110111100001110111011111111011001100111011101110111011101000111011011110111011101110100010001010111011001100110111101011111011100111111011011110100011100001111100110001111011011101110111011010011011000101111101111111101010011110111010011011011111111101011011010110001011011100111111111001111111011101101101110111111111111101111111101111111011101100111111100110000111101101111011111101101111111101111101110011001111111110011000100110111000100011111111111111100011111110001001111110111000100011111011111100111";cor_in <= "10011110101010111001100110011110010010101000000010101011101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "11111110010011000011111111111111001111111110011100111110110110000001111111111111111110001100111001110001100010000111111111111111011111111001110111111110001111111100100000011111100011001110111101110111110000001111111101110111111111111111111111111111111100011100100000001110100011111111111111111111111101101101100011111111011011111111101111111110111111111111111110000000111111111001111100111111110110011111100100111011111100000000100111110000010011001111111111110111110111111111011111111000111101111111111110110011";cor_in <= "11010100101010111001100110011110101101011000000001000000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00110111001000011111111111001111011011100100010101110110011100100111011011111111111101111101101101110111010101010011100111111111011101110110101111111111011110001111010011001011111011101000111111110111011101001001101111101110000011011111100000011111111111011111111001110111111111101111111111001111101111001111111111111111111101001100110001111011111111011111110110001000110111111111111111100111011110111011110111111111111100110100001111111111111110110111111110011100111011011111110011111111110011001001111111001101";cor_in <= "10011110101010111001100110011100010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111000011100111111111000111110011011110011011101111111111111110111111011111100111101110111011101111111011111111101011110010011111101110111110111110111111111111111110111111101110011001110111001110111111101111111001110111001100001111110000001111111110110111111101110111111111000100111111011101100110100110011111101110111011101100111010001110011101100011111111110111111111101101111011001111001011110011011101110011011111111111111111111101111111101111010011011010111001111111111000111011111110110111100111111010111";cor_in <= "10111011101010111001100101011010101101011000000010111011101000001001011110100011" ; wait for 10 ns; 
inp_feat <= "11111111100011110011110010111111000111101000001111111111111011001000111111111001111110001111111101111101111011111111111011011111111111101101111111111111111111111100111011111111100010001001001111111111111111111111111101110111110100110011011101111111111100011110111011001111110010001111100101110111001000011111111101111111000010011111100111111111111101111011100011101100101111111111011100111111110011111101111111110010111111101110011011111110110111111111100111111110100101111111000111110000111111111111100110000000";cor_in <= "01001100101010111011001010011110101111011000000010101011101000001000110110100101" ; wait for 10 ns; 
inp_feat <= "01101100010011110011111011101111011111101100000000000111111111110111111100111100011011111111011100000000111111111111111011111011011011001111011111101111101111111111111111111111111011101100000000100001111111111110110100111011110011000000000010101111000011001111111111111111111111001111000010111100000001111100000011111111011011111111000011111110001101111010111111110011111111111100011101110111000011111111111101111111101111111111111111111111111111111110100011110111110110100011000011111111011101111110110011000001";cor_in <= "10011110101010111001110010011110101111011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11111000110001100111110111111111001111111101001101101110111011100111111111101100111010001101111101110000100011110101110010001111111110001000111011111101110111011100111011111011110011001101111101110000011011101111011101100001111100110011011111111111111000111110111000000001100110011101111110111111111100011111011000101111000111011111111111111110010000001111110111111110111111011111110011111110110001110010111111110111111111001101110011111110100010011111100110111111101100110111001011110000111111111011111111010001";cor_in <= "01001100101010111010110010011100110001001001000010101011100111111000110110100101" ; wait for 10 ns; 
inp_feat <= "11110111010001010111010011011100011011111111110011110111111111111111111111111110011111101111111111110011100011111111111111111111011111111000111111111111101101110110111111111011011011001100101011110111000111111011110000110001111111110000001110111111111100011110111111111011010111001110111111111111100000001111111100111111011011001111111111111111111100111111110011111111111111111111100011111111111111011000111111110111010011111111111111111111011111111111110001001111110110100111011110101000011101111100111111111011";cor_in <= "10100010101010110100000110011110101101011000000010101011101000001000110110101011" ; wait for 10 ns; 
inp_feat <= "00110110111001100011011111101110001101110111010100000011011111001111001100101111001101101100011000000111011111100111111011110111001101101111111101111111010011111111011111001101011111111110111100010011011101101111110110010011011011101111011111111011001111000101111110001011111111101110101111011000001100111110010100110110001101111111011111001011001100111011111111111100011111011011111110110110011111101111111110110001111111111111100111011111111111000100111101100110111011000111011111111111101100011101111111110000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001010110101000000" ; wait for 10 ns; 
inp_feat <= "01000000000000001111111111101111001101100110001000100010000010101010101110101011001001100000001000000001001101110011011001110011001100000000001001100000000001101001111111001111010011000100011001100000000000001111110110011111011000000110010011101110111011101011000100010001011101110011111111101110111011101110101011101000111011101110111111111000100000000110011001100110111111111111111110111001110101111111111111111011111101110011001111010011111100010110001000100110011001100110011111111111101110110110011001100110";cor_in <= "10100010010001101001100111001101101101011000000010101011101000001000110111100000" ; wait for 10 ns; 
inp_feat <= "00001111101111111111111100111111001111100111011010111111111111111111111111111111111011110111111111111111011111110111111111111100011001110111111111101111011111111111101110011111111011001110110001111111111101111101111110011011110011001100100011010111100001110011100111111111111101111111110011001110110001111111111111111111111100110111010011101111110101111111001111110001111101111100111110001111100111111111101111111111111100111111011110101110111111111111111011111111111101111111001011111111101110111011111001110100";cor_in <= "10011110101010111001100111000001101101011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11110110111101101111110000001110011011100001011111111111111101110111111011111111111111111111011111111111111111011101111111111111111111110011010111110110111111001111111111111101110011000010111001111111111100111111001110111001100100111111111101111011111111011111111111111111110011001110111000111100111110100111011111110111111011100010111111111111111111111111111000111110111101001111110011111111111111111111011110111011111111110111111111011111111000111110011001110111001101111111011101000111011100111100111101100111";cor_in <= "10011110101010111011101101011010101101011000000010101011101000001000110110011000" ; wait for 10 ns; 
inp_feat <= "11111111011011111000000011111110100111111110100111001110011111100011111110001101111101101111111111110000111111111111111111001111111101101101011111111111111111110010011111111111000001101110100111111110011111111111111110011001111111101001001100111110000110111001111111111111000111111111111111111111001010011111101100111111000000101111110011111111111100111110000111110000011111111110001111111111111011110011111111011011101111111111001111111101011111111110000101110110111111110011000111110011011101111110110111010000";cor_in <= "10011110101010110100010010011110101101011000000010101011101001111000110110000001" ; wait for 10 ns; 
inp_feat <= "00000011111101110011011111101110011101110111011101110011111011001111101101111111011111101110111000100111001111001111111110111111001001111111111001111110111100111111011110101101001111111111111101100011011101001101110110111010011011011111011011111011001111100101111111011111111111111111111011101100111100111110111100110101011101111111000011101111111100111011111011001100111101101111111111111001111111111111111100010001111111111001100110001110111011110110111111110100111111110111001111011111101100111111001101100110";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 
inp_feat <= "00110000100111110001011111001111001101111110110100000011111111111011011100001110011111111111111100110011011111111111111001110110001000001011111111111111111111111111111111001111011111101110111000110001011101111101111100010111111011101111000011111001000101101101101101111111111111101110100011011010101000111111111101111111001101111111000011111111001111111111111111110001111110011011011110110111000111111101111110110011100111111111011111111111111111111101110011111111111111111011000011111111111101111011100011110000";cor_in <= "11000010101010111001100110011110110011011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "00110001000011101100111111111111111111110111001100110101111011100111011001011111010101011111111011010100111111110110111101111111000000110111011100110111011111101111110110101111011001100101011111010011111111101011111110011010010000001011000011011111011111110011001100001111011011100111110111111111111110111011100111111111111011111111010101111111000101111111001111110000111111111111111111111101101111111111111111111111111111111111000100110011000001000100011111100111111111101111000111110111111111011111111101110001";cor_in <= "10011110101010111001100110011110101101011000000010101011001110011000110110101000" ; wait for 10 ns; 
inp_feat <= "11111110100000100011111110110011001101111111111111111111110001000000111111111011111111001100011001111111110000000111011111111111111111010100001011110011011011010000110011101111110011100101011101111110000000001111011101111101111111110111011001111111111111111100100011001101110010110011111111110111011111010110110111101111111011110011001111110110111111101111111100001110111110110011110101111111111010110011000111111111111000011001110011111001110011101111011100111110110101111111111111111101001111111111011111011110";cor_in <= "10011110101010111001100110011110101101011000100001000000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111000000011001001111111100000001111111110011101111011101110000111111110110111101110001111111111111000011111101111111111111111101110000111111110111111101100000011111111001001001111100111011111000000001111101111111000011111111101100001000011110111100010110111111110111001100001110111011011111100010001111111110110111001100001111111100011111111111111111000111011111111111011111110010111111111110011101001111111011111100011111111111111111011101111111110011000111110111010111111111111001000101111011110011111111";cor_in <= "10011110101010110100010010011110101101011000000010101011101000001000110110111100" ; wait for 10 ns; 
inp_feat <= "00000000000111111110110011111111111011110110110100000111011111100111011101101100000001011111111100000000111111110110111011111111000000000111011101100111111111111101110111111111111010001111110100000000011111111011101110010010110011011101001011111101011111110011001101111111011111101111110011001111111001111011111101111111111011101111110101001111111100110111011111110001111111111111101100110111100111111111111111111110011111111111001100110011000111011100111111110100110111111110000010111111111111111101111101110101";cor_in <= "10011110101010111001100110011110101101011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11001111011111111111111100001101011110110010011111111111111011001011110111111111110111111111111111111111001100111011111111111111111101110111111111111110111111111000111100001111110010111110111101111111111100100111001011110111001111101111111111111101111100111100000110001111111110111111111111101101101101110100110101111011111110110111110011111110111111111111101110011100111100110000100111111111111111110011110111011000101100111001000000011111111111110111111111111110011111111111001111010101001111101111001100000000";cor_in <= "10011110101010111001100110011110101101011000000010101011101000000011111110000001" ; wait for 10 ns; 
inp_feat <= "10000011011100001111110000011111011011111111111101110001011001100111100011110111111111111110100001110111011101011110100110001111010101110111110111110111111010110111100011101111111011101111110011011111001101001111000111111110110011011111111011011001111111111011111111111110111111111101111011001101111111111111111100100010111101110101110111110001011101111111111100111101111011111111100111101001011111111011101111001100011111110011100010111111111101001011011100010101111111001011000011111111111000001101111111011101";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00000000000011111111011111111111001101100111110000000011011111111011011100111110011001111111111100010010011111110111111010111001000000001111011101101111011111111111011111111111001111101110110000000000011111111111111110010001111011001000000011111111000111011001101111111111111111101110100011111111100001111100110101111111011101100111000010100001001101111111011111110011011111111110011111010111000111111111111110111001101111111111111111011100011111111100110011110111111011001110000111111111111111111111110001110111";cor_in <= "10011110101010111001100110011110101101011000000010101011010001011000110110000001" ; wait for 10 ns; 
inp_feat <= "11110110111100111111111110011111011111101111001111111111111111111111101111111110111111110011011111101111111101111111111111111111111111011111011111111111111101111101111110111110111011101001011101110111111111110011000110011101111010010111111011110001101111001111111110111111111111100111111100100110111110000110011111110011111011110011101111111111101111011111111100110011111111101111111001111110111111011001011110011001111111110011111111010111111110111110111101110011101100111111011111110111001100111100111101100011";cor_in <= "10011110101010111001100101011010101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111110000000001100111110111101111110111111111111111100011001000111111011101111110001100001001110111110100000111111111101111111111111101000111101111011101010001000011101111110011101110001101111110101010101111011101101111111101111011101110111111011111111000110011001100100011111111011111111111111101101110110111111110111111110111001111111111011011111111101100010100111110111111111101111111111011001111000111111111111000010001110111111101110011001111111100110011110111110111111111110001011111111111101100111111";cor_in <= "10011110101010111001100110011110101101011000011001000000101011001000110110000001" ; wait for 10 ns; 
inp_feat <= "00000000000000000111111110001110111111111110111000000000000001101011100111110011001100100100110000110000001000001101011110101110001100000010010001110110011011001110111111111111000011111110111001100000000000101111111111111011011101101100110011111110111011100111111110111111011111111111111011101100111111100010111111001110011111110010111010111000010101101111011001101100111111110111111110111011001011101011111111111111111111111011111111111111111101110110011011101110011101111110100011111111111100110110111111100110";cor_in <= "10111110010001101001100110011110101101011001011110101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11100100111111110111111110001100011011101101011101110111111111110111011101111111110111111111111100111111111110111101111111111111111111100111111111110110111111111111111100011100110011000010111001110111111111111111001110110011111100001111101101110111101110111110111100111111110011101110111010111000111000110111011101110111111111111111010011111111011110111111111011101110111111011110110101111111111111111111111100110011110011110111110111001111111111111111111111111110101111111111011111001111111101111100111111000111";cor_in <= "10011110101010111001110001011010101101011000000010101011101000001001000010010001" ; wait for 10 ns; 
inp_feat <= "11111111110000000011110111000001001101110111011101111110111011000000111111111111111011001100111001111111110000001111111111111111111111111111001011101111011111100000100011101111100011101111011111110111111000001111001101111111111101111111111010111111111111111100110001101111100011110111111111101111011111110111011011101110011111110001011111110111011111111111110100001000111110110011111111111111111110000111000111011111111111011001100111110111111011101111011101111111111101110111111111110101000101111111001100101110";cor_in <= "10011110101010111001100110011110101101011010011001000000101001111000110110100101" ; wait for 10 ns; 
inp_feat <= "00110111011111000011101101001110001100111111111101110011111011001011010011111111111101111100110000110011001001000111111111111111001101111111111001111100111110001111110111001111011101101111111100010011001101101101101111011011011011011111111000110011111000101111111011111111011111101111111111001111011100111111101100110100011101111111111011111111111111111111111110001100011111101011001110011011111111111111111111010101111111011001100111101110111011110111111111111100111111111111111111111111101101110001011110000000";cor_in <= "10011110101010111001100110011110101111011000000010101011101000001000110100011110" ; wait for 10 ns; 
inp_feat <= "11110000011101111111111011111111011011110101001101110111110111010111011110111111011101100111011100110111111111111101011110111001011100010111111111110110111101101111111110001111111011001000111101110011111101111111101110111001110100001011001011110111100110011111111110011111110011000111101111101100110000100111001100110111011001100111011101110111001100010111111011110111111111111111011001111111101110011011101110010001111111111111111111111111111110111110011011101111010001011101001111011111110110011100111111100011";cor_in <= "10011011101010111001100101011010101101011000000010101011101000001000110110110000" ; wait for 10 ns; 
inp_feat <= "11100000000000001110101110111111011100110111011110000000000011101000101111111011010000000000010011110110011101110011100110111001011000000000001011101100010001101000110011001100000001110111010011110100000001111111111110011101011001100100011011111110101011111010100110011101011101111111101111001110111011100110100010001001011011111111111101110000000000001111011001100111111101111111111110111011111111111111111111111011111111111101011111111010001100111110101000100010010101100110011110111101101110111110111001110111";cor_in <= "10011110010001101001100110011110101101011001000110101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "11111111110011101111000111001110001101101111111111111110111111001011011111111111111110011100111001110111001100001011110001111111011111111111111111111111110111111101000010011111000011101111111111111111001110001011110111110101111011111111111010011101101011011011100010001111111111000111111111001011111100110111111110101011011100010101100001110101111110111111111111000000111110110001100110111111111111111101100100010001111110010000000111111111101010111001111101111110111011111111111111111111000010011101101100001001";cor_in <= "10011110101010111001100110011110010110011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "01100010001100011110111111101111011011100111000101100010111111111110101110101111111011100110000011101111111111110010011001111001011001100110001110100100010001001001100111011110110001100110000011100110011111111111101110011101000001000000001011111011111111010011000110011000011001100111011111001110111011100100100010001010111011111111111111000000000000011111111101110011111101111111101111101111110101111111101111111001111101110111101000010001100110010110001001100011111011110111011111111011101110111110111001100011";cor_in <= "10011110110100101001100110011110101101011000000010101011101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00001101111111111111011100011111001101111111011111111001111111111111001111111100111011111111111111111111111101110011111111101111000011101111011111101110111111111101000110111111001111110110111011101111111100111111110111011001011011101110110111111101100110110001100111111111111101110011111011101100111100111100110111111011111111110111011011001100110111111111111001110111111101101111011111110011111111011111110110111001111110001111100110011011111101110000111100111111111011111111000011011111000110110111001101010111";cor_in <= "10011110101010111001100110011110101101011000000010101011010001011100001010000001" ; wait for 10 ns; 
inp_feat <= "11111110000010001101110101011111001101111111001111111110110011001110111111111011111111001110111011111111100011000011111111110111111111110001111111101011111111001000110011111111110010100001111111111111110011100011011111111111111111111111011000111111111101101100111011101001110010010001111101110111011110110110111111101111111100010011111111110111111111111111000110001100101100111111100111111111111011110011110111111111110011011100100011111110110011001111001101111111011100111111111111110000111111110111001111111001";cor_in <= "10011110101010111001100110011110101111001000000001000000101000001000110110000001" ; wait for 10 ns; 
inp_feat <= "00111111111011111111110111111111011101111110100101110011011011100111010011111111111111111100011111110111111111110111111110111111001100111110011101111111111011111111000011001111011011101111011110110111001111111011101100111001110011110011001111010111011110010011111010101101011011001111101111001011011100111011111100110110111111100111010111111111011100111111111111110100111111111111010011000111111111111111101110011000111110111100100111111111011011111111111101100110111011110011000111111111010000111111011111000001";cor_in <= "10011110101010111001100110011110101101011000000010101011101000001000110101000000" ; wait for 10 ns; 

      -- insert stimulus here 

      wait;
   end process;

END;
