----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:45:07 07/27/2019 
-- Design Name: 
-- Module Name:    SVHN_full_check - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity svhn_reg_fin is
    Port ( inp_feat : in  STD_LOGIC_VECTOR (511 downto 0);
           out_fin : out  STD_LOGIC_VECTOR (79 downto 0));
           --cor_in : in  STD_LOGIC_VECTOR (79 downto 0);
           --cor_out : out  STD_LOGIC_VECTOR (79 downto 0));
end svhn_reg_fin;

architecture Behavioral of svhn_reg_fin is

signal C_0_out : std_logic := '0'; 
signal C_1_out : std_logic := '0'; 
signal C_2_out : std_logic := '0'; 
signal C_3_out : std_logic := '0'; 
signal C_4_out : std_logic := '0'; 
signal C_5_out : std_logic := '0'; 
signal C_6_out : std_logic := '0'; 
signal C_7_out : std_logic := '0'; 
signal C_8_out : std_logic := '0'; 
signal C_9_out : std_logic := '0'; 
signal C_10_out : std_logic := '0'; 
signal C_11_out : std_logic := '0'; 
signal C_12_out : std_logic := '0'; 
signal C_13_out : std_logic := '0'; 
signal C_14_out : std_logic := '0'; 
signal C_15_out : std_logic := '0'; 
signal C_16_out : std_logic := '0'; 
signal C_17_out : std_logic := '0'; 
signal C_18_out : std_logic := '0'; 
signal C_19_out : std_logic := '0'; 
signal C_20_out : std_logic := '0'; 
signal C_21_out : std_logic := '0'; 
signal C_22_out : std_logic := '0'; 
signal C_23_out : std_logic := '0'; 
signal C_24_out : std_logic := '0'; 
signal C_25_out : std_logic := '0'; 
signal C_26_out : std_logic := '0'; 
signal C_27_out : std_logic := '0'; 
signal C_28_out : std_logic := '0'; 
signal C_29_out : std_logic := '0'; 
signal C_30_out : std_logic := '0'; 
signal C_31_out : std_logic := '0'; 
signal C_32_out : std_logic := '0'; 
signal C_33_out : std_logic := '0'; 
signal C_34_out : std_logic := '0'; 
signal C_35_out : std_logic := '0'; 
signal C_36_out : std_logic := '0'; 
signal C_37_out : std_logic := '0'; 
signal C_38_out : std_logic := '0'; 
signal C_39_out : std_logic := '0'; 
signal C_40_out : std_logic := '0'; 
signal C_41_out : std_logic := '0'; 
signal C_42_out : std_logic := '0'; 
signal C_43_out : std_logic := '0'; 
signal C_44_out : std_logic := '0'; 
signal C_45_out : std_logic := '0'; 
signal C_46_out : std_logic := '0'; 
signal C_47_out : std_logic := '0'; 
signal C_48_out : std_logic := '0'; 
signal C_49_out : std_logic := '0'; 
signal C_50_out : std_logic := '0'; 
signal C_51_out : std_logic := '0'; 
signal C_52_out : std_logic := '0'; 
signal C_53_out : std_logic := '0'; 
signal C_54_out : std_logic := '0'; 
signal C_55_out : std_logic := '0'; 
signal C_56_out : std_logic := '0'; 
signal C_57_out : std_logic := '0'; 
signal C_58_out : std_logic := '0'; 
signal C_59_out : std_logic := '0'; 

signal C_0_S_0_L_0_out : std_logic := '0'; 
signal C_0_S_0_L_1_out : std_logic := '0'; 
signal C_0_S_0_L_2_out : std_logic := '0'; 
signal C_0_S_0_L_3_out : std_logic := '0'; 
signal C_0_S_0_L_4_out : std_logic := '0'; 
signal C_0_S_0_L_5_out : std_logic := '0'; 
signal C_0_S_1_L_0_out : std_logic := '0'; 
signal C_0_S_1_L_1_out : std_logic := '0'; 
signal C_0_S_1_L_2_out : std_logic := '0'; 
signal C_0_S_1_L_3_out : std_logic := '0'; 
signal C_0_S_1_L_4_out : std_logic := '0'; 
signal C_0_S_1_L_5_out : std_logic := '0'; 
signal C_0_S_2_L_0_out : std_logic := '0'; 
signal C_0_S_2_L_1_out : std_logic := '0'; 
signal C_0_S_2_L_2_out : std_logic := '0'; 
signal C_0_S_2_L_3_out : std_logic := '0'; 
signal C_0_S_2_L_4_out : std_logic := '0'; 
signal C_0_S_2_L_5_out : std_logic := '0'; 
signal C_0_S_3_L_0_out : std_logic := '0'; 
signal C_0_S_3_L_1_out : std_logic := '0'; 
signal C_0_S_3_L_2_out : std_logic := '0'; 
signal C_0_S_3_L_3_out : std_logic := '0'; 
signal C_0_S_3_L_4_out : std_logic := '0'; 
signal C_0_S_3_L_5_out : std_logic := '0'; 
signal C_0_S_4_L_0_out : std_logic := '0'; 
signal C_0_S_4_L_1_out : std_logic := '0'; 
signal C_0_S_4_L_2_out : std_logic := '0'; 
signal C_0_S_4_L_3_out : std_logic := '0'; 
signal C_0_S_4_L_4_out : std_logic := '0'; 
signal C_0_S_4_L_5_out : std_logic := '0'; 
signal C_0_S_5_L_0_out : std_logic := '0'; 
signal C_0_S_5_L_1_out : std_logic := '0'; 
signal C_0_S_5_L_2_out : std_logic := '0'; 
signal C_0_S_5_L_3_out : std_logic := '0'; 
signal C_0_S_5_L_4_out : std_logic := '0'; 
signal C_0_S_5_L_5_out : std_logic := '0'; 
signal C_1_S_0_L_0_out : std_logic := '0'; 
signal C_1_S_0_L_1_out : std_logic := '0'; 
signal C_1_S_0_L_2_out : std_logic := '0'; 
signal C_1_S_0_L_3_out : std_logic := '0'; 
signal C_1_S_0_L_4_out : std_logic := '0'; 
signal C_1_S_0_L_5_out : std_logic := '0'; 
signal C_1_S_1_L_0_out : std_logic := '0'; 
signal C_1_S_1_L_1_out : std_logic := '0'; 
signal C_1_S_1_L_2_out : std_logic := '0'; 
signal C_1_S_1_L_3_out : std_logic := '0'; 
signal C_1_S_1_L_4_out : std_logic := '0'; 
signal C_1_S_1_L_5_out : std_logic := '0'; 
signal C_1_S_2_L_0_out : std_logic := '0'; 
signal C_1_S_2_L_1_out : std_logic := '0'; 
signal C_1_S_2_L_2_out : std_logic := '0'; 
signal C_1_S_2_L_3_out : std_logic := '0'; 
signal C_1_S_2_L_4_out : std_logic := '0'; 
signal C_1_S_2_L_5_out : std_logic := '0'; 
signal C_1_S_3_L_0_out : std_logic := '0'; 
signal C_1_S_3_L_1_out : std_logic := '0'; 
signal C_1_S_3_L_2_out : std_logic := '0'; 
signal C_1_S_3_L_3_out : std_logic := '0'; 
signal C_1_S_3_L_4_out : std_logic := '0'; 
signal C_1_S_3_L_5_out : std_logic := '0'; 
signal C_1_S_4_L_0_out : std_logic := '0'; 
signal C_1_S_4_L_1_out : std_logic := '0'; 
signal C_1_S_4_L_2_out : std_logic := '0'; 
signal C_1_S_4_L_3_out : std_logic := '0'; 
signal C_1_S_4_L_4_out : std_logic := '0'; 
signal C_1_S_4_L_5_out : std_logic := '0'; 
signal C_1_S_5_L_0_out : std_logic := '0'; 
signal C_1_S_5_L_1_out : std_logic := '0'; 
signal C_1_S_5_L_2_out : std_logic := '0'; 
signal C_1_S_5_L_3_out : std_logic := '0'; 
signal C_1_S_5_L_4_out : std_logic := '0'; 
signal C_1_S_5_L_5_out : std_logic := '0'; 
signal C_2_S_0_L_0_out : std_logic := '0'; 
signal C_2_S_0_L_1_out : std_logic := '0'; 
signal C_2_S_0_L_2_out : std_logic := '0'; 
signal C_2_S_0_L_3_out : std_logic := '0'; 
signal C_2_S_0_L_4_out : std_logic := '0'; 
signal C_2_S_0_L_5_out : std_logic := '0'; 
signal C_2_S_1_L_0_out : std_logic := '0'; 
signal C_2_S_1_L_1_out : std_logic := '0'; 
signal C_2_S_1_L_2_out : std_logic := '0'; 
signal C_2_S_1_L_3_out : std_logic := '0'; 
signal C_2_S_1_L_4_out : std_logic := '0'; 
signal C_2_S_1_L_5_out : std_logic := '0'; 
signal C_2_S_2_L_0_out : std_logic := '0'; 
signal C_2_S_2_L_1_out : std_logic := '0'; 
signal C_2_S_2_L_2_out : std_logic := '0'; 
signal C_2_S_2_L_3_out : std_logic := '0'; 
signal C_2_S_2_L_4_out : std_logic := '0'; 
signal C_2_S_2_L_5_out : std_logic := '0'; 
signal C_2_S_3_L_0_out : std_logic := '0'; 
signal C_2_S_3_L_1_out : std_logic := '0'; 
signal C_2_S_3_L_2_out : std_logic := '0'; 
signal C_2_S_3_L_3_out : std_logic := '0'; 
signal C_2_S_3_L_4_out : std_logic := '0'; 
signal C_2_S_3_L_5_out : std_logic := '0'; 
signal C_2_S_4_L_0_out : std_logic := '0'; 
signal C_2_S_4_L_1_out : std_logic := '0'; 
signal C_2_S_4_L_2_out : std_logic := '0'; 
signal C_2_S_4_L_3_out : std_logic := '0'; 
signal C_2_S_4_L_4_out : std_logic := '0'; 
signal C_2_S_4_L_5_out : std_logic := '0'; 
signal C_2_S_5_L_0_out : std_logic := '0'; 
signal C_2_S_5_L_1_out : std_logic := '0'; 
signal C_2_S_5_L_2_out : std_logic := '0'; 
signal C_2_S_5_L_3_out : std_logic := '0'; 
signal C_2_S_5_L_4_out : std_logic := '0'; 
signal C_2_S_5_L_5_out : std_logic := '0'; 
signal C_3_S_0_L_0_out : std_logic := '0'; 
signal C_3_S_0_L_1_out : std_logic := '0'; 
signal C_3_S_0_L_2_out : std_logic := '0'; 
signal C_3_S_0_L_3_out : std_logic := '0'; 
signal C_3_S_0_L_4_out : std_logic := '0'; 
signal C_3_S_0_L_5_out : std_logic := '0'; 
signal C_3_S_1_L_0_out : std_logic := '0'; 
signal C_3_S_1_L_1_out : std_logic := '0'; 
signal C_3_S_1_L_2_out : std_logic := '0'; 
signal C_3_S_1_L_3_out : std_logic := '0'; 
signal C_3_S_1_L_4_out : std_logic := '0'; 
signal C_3_S_1_L_5_out : std_logic := '0'; 
signal C_3_S_2_L_0_out : std_logic := '0'; 
signal C_3_S_2_L_1_out : std_logic := '0'; 
signal C_3_S_2_L_2_out : std_logic := '0'; 
signal C_3_S_2_L_3_out : std_logic := '0'; 
signal C_3_S_2_L_4_out : std_logic := '0'; 
signal C_3_S_2_L_5_out : std_logic := '0'; 
signal C_3_S_3_L_0_out : std_logic := '0'; 
signal C_3_S_3_L_1_out : std_logic := '0'; 
signal C_3_S_3_L_2_out : std_logic := '0'; 
signal C_3_S_3_L_3_out : std_logic := '0'; 
signal C_3_S_3_L_4_out : std_logic := '0'; 
signal C_3_S_3_L_5_out : std_logic := '0'; 
signal C_3_S_4_L_0_out : std_logic := '0'; 
signal C_3_S_4_L_1_out : std_logic := '0'; 
signal C_3_S_4_L_2_out : std_logic := '0'; 
signal C_3_S_4_L_3_out : std_logic := '0'; 
signal C_3_S_4_L_4_out : std_logic := '0'; 
signal C_3_S_4_L_5_out : std_logic := '0'; 
signal C_3_S_5_L_0_out : std_logic := '0'; 
signal C_3_S_5_L_1_out : std_logic := '0'; 
signal C_3_S_5_L_2_out : std_logic := '0'; 
signal C_3_S_5_L_3_out : std_logic := '0'; 
signal C_3_S_5_L_4_out : std_logic := '0'; 
signal C_3_S_5_L_5_out : std_logic := '0'; 
signal C_4_S_0_L_0_out : std_logic := '0'; 
signal C_4_S_0_L_1_out : std_logic := '0'; 
signal C_4_S_0_L_2_out : std_logic := '0'; 
signal C_4_S_0_L_3_out : std_logic := '0'; 
signal C_4_S_0_L_4_out : std_logic := '0'; 
signal C_4_S_0_L_5_out : std_logic := '0'; 
signal C_4_S_1_L_0_out : std_logic := '0'; 
signal C_4_S_1_L_1_out : std_logic := '0'; 
signal C_4_S_1_L_2_out : std_logic := '0'; 
signal C_4_S_1_L_3_out : std_logic := '0'; 
signal C_4_S_1_L_4_out : std_logic := '0'; 
signal C_4_S_1_L_5_out : std_logic := '0'; 
signal C_4_S_2_L_0_out : std_logic := '0'; 
signal C_4_S_2_L_1_out : std_logic := '0'; 
signal C_4_S_2_L_2_out : std_logic := '0'; 
signal C_4_S_2_L_3_out : std_logic := '0'; 
signal C_4_S_2_L_4_out : std_logic := '0'; 
signal C_4_S_2_L_5_out : std_logic := '0'; 
signal C_4_S_3_L_0_out : std_logic := '0'; 
signal C_4_S_3_L_1_out : std_logic := '0'; 
signal C_4_S_3_L_2_out : std_logic := '0'; 
signal C_4_S_3_L_3_out : std_logic := '0'; 
signal C_4_S_3_L_4_out : std_logic := '0'; 
signal C_4_S_3_L_5_out : std_logic := '0'; 
signal C_4_S_4_L_0_out : std_logic := '0'; 
signal C_4_S_4_L_1_out : std_logic := '0'; 
signal C_4_S_4_L_2_out : std_logic := '0'; 
signal C_4_S_4_L_3_out : std_logic := '0'; 
signal C_4_S_4_L_4_out : std_logic := '0'; 
signal C_4_S_4_L_5_out : std_logic := '0'; 
signal C_4_S_5_L_0_out : std_logic := '0'; 
signal C_4_S_5_L_1_out : std_logic := '0'; 
signal C_4_S_5_L_2_out : std_logic := '0'; 
signal C_4_S_5_L_3_out : std_logic := '0'; 
signal C_4_S_5_L_4_out : std_logic := '0'; 
signal C_4_S_5_L_5_out : std_logic := '0'; 
signal C_5_S_0_L_0_out : std_logic := '0'; 
signal C_5_S_0_L_1_out : std_logic := '0'; 
signal C_5_S_0_L_2_out : std_logic := '0'; 
signal C_5_S_0_L_3_out : std_logic := '0'; 
signal C_5_S_0_L_4_out : std_logic := '0'; 
signal C_5_S_0_L_5_out : std_logic := '0'; 
signal C_5_S_1_L_0_out : std_logic := '0'; 
signal C_5_S_1_L_1_out : std_logic := '0'; 
signal C_5_S_1_L_2_out : std_logic := '0'; 
signal C_5_S_1_L_3_out : std_logic := '0'; 
signal C_5_S_1_L_4_out : std_logic := '0'; 
signal C_5_S_1_L_5_out : std_logic := '0'; 
signal C_5_S_2_L_0_out : std_logic := '0'; 
signal C_5_S_2_L_1_out : std_logic := '0'; 
signal C_5_S_2_L_2_out : std_logic := '0'; 
signal C_5_S_2_L_3_out : std_logic := '0'; 
signal C_5_S_2_L_4_out : std_logic := '0'; 
signal C_5_S_2_L_5_out : std_logic := '0'; 
signal C_5_S_3_L_0_out : std_logic := '0'; 
signal C_5_S_3_L_1_out : std_logic := '0'; 
signal C_5_S_3_L_2_out : std_logic := '0'; 
signal C_5_S_3_L_3_out : std_logic := '0'; 
signal C_5_S_3_L_4_out : std_logic := '0'; 
signal C_5_S_3_L_5_out : std_logic := '0'; 
signal C_5_S_4_L_0_out : std_logic := '0'; 
signal C_5_S_4_L_1_out : std_logic := '0'; 
signal C_5_S_4_L_2_out : std_logic := '0'; 
signal C_5_S_4_L_3_out : std_logic := '0'; 
signal C_5_S_4_L_4_out : std_logic := '0'; 
signal C_5_S_4_L_5_out : std_logic := '0'; 
signal C_5_S_5_L_0_out : std_logic := '0'; 
signal C_5_S_5_L_1_out : std_logic := '0'; 
signal C_5_S_5_L_2_out : std_logic := '0'; 
signal C_5_S_5_L_3_out : std_logic := '0'; 
signal C_5_S_5_L_4_out : std_logic := '0'; 
signal C_5_S_5_L_5_out : std_logic := '0'; 
signal C_6_S_0_L_0_out : std_logic := '0'; 
signal C_6_S_0_L_1_out : std_logic := '0'; 
signal C_6_S_0_L_2_out : std_logic := '0'; 
signal C_6_S_0_L_3_out : std_logic := '0'; 
signal C_6_S_0_L_4_out : std_logic := '0'; 
signal C_6_S_0_L_5_out : std_logic := '0'; 
signal C_6_S_1_L_0_out : std_logic := '0'; 
signal C_6_S_1_L_1_out : std_logic := '0'; 
signal C_6_S_1_L_2_out : std_logic := '0'; 
signal C_6_S_1_L_3_out : std_logic := '0'; 
signal C_6_S_1_L_4_out : std_logic := '0'; 
signal C_6_S_1_L_5_out : std_logic := '0'; 
signal C_6_S_2_L_0_out : std_logic := '0'; 
signal C_6_S_2_L_1_out : std_logic := '0'; 
signal C_6_S_2_L_2_out : std_logic := '0'; 
signal C_6_S_2_L_3_out : std_logic := '0'; 
signal C_6_S_2_L_4_out : std_logic := '0'; 
signal C_6_S_2_L_5_out : std_logic := '0'; 
signal C_6_S_3_L_0_out : std_logic := '0'; 
signal C_6_S_3_L_1_out : std_logic := '0'; 
signal C_6_S_3_L_2_out : std_logic := '0'; 
signal C_6_S_3_L_3_out : std_logic := '0'; 
signal C_6_S_3_L_4_out : std_logic := '0'; 
signal C_6_S_3_L_5_out : std_logic := '0'; 
signal C_6_S_4_L_0_out : std_logic := '0'; 
signal C_6_S_4_L_1_out : std_logic := '0'; 
signal C_6_S_4_L_2_out : std_logic := '0'; 
signal C_6_S_4_L_3_out : std_logic := '0'; 
signal C_6_S_4_L_4_out : std_logic := '0'; 
signal C_6_S_4_L_5_out : std_logic := '0'; 
signal C_6_S_5_L_0_out : std_logic := '0'; 
signal C_6_S_5_L_1_out : std_logic := '0'; 
signal C_6_S_5_L_2_out : std_logic := '0'; 
signal C_6_S_5_L_3_out : std_logic := '0'; 
signal C_6_S_5_L_4_out : std_logic := '0'; 
signal C_6_S_5_L_5_out : std_logic := '0'; 
signal C_7_S_0_L_0_out : std_logic := '0'; 
signal C_7_S_0_L_1_out : std_logic := '0'; 
signal C_7_S_0_L_2_out : std_logic := '0'; 
signal C_7_S_0_L_3_out : std_logic := '0'; 
signal C_7_S_0_L_4_out : std_logic := '0'; 
signal C_7_S_0_L_5_out : std_logic := '0'; 
signal C_7_S_1_L_0_out : std_logic := '0'; 
signal C_7_S_1_L_1_out : std_logic := '0'; 
signal C_7_S_1_L_2_out : std_logic := '0'; 
signal C_7_S_1_L_3_out : std_logic := '0'; 
signal C_7_S_1_L_4_out : std_logic := '0'; 
signal C_7_S_1_L_5_out : std_logic := '0'; 
signal C_7_S_2_L_0_out : std_logic := '0'; 
signal C_7_S_2_L_1_out : std_logic := '0'; 
signal C_7_S_2_L_2_out : std_logic := '0'; 
signal C_7_S_2_L_3_out : std_logic := '0'; 
signal C_7_S_2_L_4_out : std_logic := '0'; 
signal C_7_S_2_L_5_out : std_logic := '0'; 
signal C_7_S_3_L_0_out : std_logic := '0'; 
signal C_7_S_3_L_1_out : std_logic := '0'; 
signal C_7_S_3_L_2_out : std_logic := '0'; 
signal C_7_S_3_L_3_out : std_logic := '0'; 
signal C_7_S_3_L_4_out : std_logic := '0'; 
signal C_7_S_3_L_5_out : std_logic := '0'; 
signal C_7_S_4_L_0_out : std_logic := '0'; 
signal C_7_S_4_L_1_out : std_logic := '0'; 
signal C_7_S_4_L_2_out : std_logic := '0'; 
signal C_7_S_4_L_3_out : std_logic := '0'; 
signal C_7_S_4_L_4_out : std_logic := '0'; 
signal C_7_S_4_L_5_out : std_logic := '0'; 
signal C_7_S_5_L_0_out : std_logic := '0'; 
signal C_7_S_5_L_1_out : std_logic := '0'; 
signal C_7_S_5_L_2_out : std_logic := '0'; 
signal C_7_S_5_L_3_out : std_logic := '0'; 
signal C_7_S_5_L_4_out : std_logic := '0'; 
signal C_7_S_5_L_5_out : std_logic := '0'; 
signal C_8_S_0_L_0_out : std_logic := '0'; 
signal C_8_S_0_L_1_out : std_logic := '0'; 
signal C_8_S_0_L_2_out : std_logic := '0'; 
signal C_8_S_0_L_3_out : std_logic := '0'; 
signal C_8_S_0_L_4_out : std_logic := '0'; 
signal C_8_S_0_L_5_out : std_logic := '0'; 
signal C_8_S_1_L_0_out : std_logic := '0'; 
signal C_8_S_1_L_1_out : std_logic := '0'; 
signal C_8_S_1_L_2_out : std_logic := '0'; 
signal C_8_S_1_L_3_out : std_logic := '0'; 
signal C_8_S_1_L_4_out : std_logic := '0'; 
signal C_8_S_1_L_5_out : std_logic := '0'; 
signal C_8_S_2_L_0_out : std_logic := '0'; 
signal C_8_S_2_L_1_out : std_logic := '0'; 
signal C_8_S_2_L_2_out : std_logic := '0'; 
signal C_8_S_2_L_3_out : std_logic := '0'; 
signal C_8_S_2_L_4_out : std_logic := '0'; 
signal C_8_S_2_L_5_out : std_logic := '0'; 
signal C_8_S_3_L_0_out : std_logic := '0'; 
signal C_8_S_3_L_1_out : std_logic := '0'; 
signal C_8_S_3_L_2_out : std_logic := '0'; 
signal C_8_S_3_L_3_out : std_logic := '0'; 
signal C_8_S_3_L_4_out : std_logic := '0'; 
signal C_8_S_3_L_5_out : std_logic := '0'; 
signal C_8_S_4_L_0_out : std_logic := '0'; 
signal C_8_S_4_L_1_out : std_logic := '0'; 
signal C_8_S_4_L_2_out : std_logic := '0'; 
signal C_8_S_4_L_3_out : std_logic := '0'; 
signal C_8_S_4_L_4_out : std_logic := '0'; 
signal C_8_S_4_L_5_out : std_logic := '0'; 
signal C_8_S_5_L_0_out : std_logic := '0'; 
signal C_8_S_5_L_1_out : std_logic := '0'; 
signal C_8_S_5_L_2_out : std_logic := '0'; 
signal C_8_S_5_L_3_out : std_logic := '0'; 
signal C_8_S_5_L_4_out : std_logic := '0'; 
signal C_8_S_5_L_5_out : std_logic := '0'; 
signal C_9_S_0_L_0_out : std_logic := '0'; 
signal C_9_S_0_L_1_out : std_logic := '0'; 
signal C_9_S_0_L_2_out : std_logic := '0'; 
signal C_9_S_0_L_3_out : std_logic := '0'; 
signal C_9_S_0_L_4_out : std_logic := '0'; 
signal C_9_S_0_L_5_out : std_logic := '0'; 
signal C_9_S_1_L_0_out : std_logic := '0'; 
signal C_9_S_1_L_1_out : std_logic := '0'; 
signal C_9_S_1_L_2_out : std_logic := '0'; 
signal C_9_S_1_L_3_out : std_logic := '0'; 
signal C_9_S_1_L_4_out : std_logic := '0'; 
signal C_9_S_1_L_5_out : std_logic := '0'; 
signal C_9_S_2_L_0_out : std_logic := '0'; 
signal C_9_S_2_L_1_out : std_logic := '0'; 
signal C_9_S_2_L_2_out : std_logic := '0'; 
signal C_9_S_2_L_3_out : std_logic := '0'; 
signal C_9_S_2_L_4_out : std_logic := '0'; 
signal C_9_S_2_L_5_out : std_logic := '0'; 
signal C_9_S_3_L_0_out : std_logic := '0'; 
signal C_9_S_3_L_1_out : std_logic := '0'; 
signal C_9_S_3_L_2_out : std_logic := '0'; 
signal C_9_S_3_L_3_out : std_logic := '0'; 
signal C_9_S_3_L_4_out : std_logic := '0'; 
signal C_9_S_3_L_5_out : std_logic := '0'; 
signal C_9_S_4_L_0_out : std_logic := '0'; 
signal C_9_S_4_L_1_out : std_logic := '0'; 
signal C_9_S_4_L_2_out : std_logic := '0'; 
signal C_9_S_4_L_3_out : std_logic := '0'; 
signal C_9_S_4_L_4_out : std_logic := '0'; 
signal C_9_S_4_L_5_out : std_logic := '0'; 
signal C_9_S_5_L_0_out : std_logic := '0'; 
signal C_9_S_5_L_1_out : std_logic := '0'; 
signal C_9_S_5_L_2_out : std_logic := '0'; 
signal C_9_S_5_L_3_out : std_logic := '0'; 
signal C_9_S_5_L_4_out : std_logic := '0'; 
signal C_9_S_5_L_5_out : std_logic := '0'; 
signal C_10_S_0_L_0_out : std_logic := '0'; 
signal C_10_S_0_L_1_out : std_logic := '0'; 
signal C_10_S_0_L_2_out : std_logic := '0'; 
signal C_10_S_0_L_3_out : std_logic := '0'; 
signal C_10_S_0_L_4_out : std_logic := '0'; 
signal C_10_S_0_L_5_out : std_logic := '0'; 
signal C_10_S_1_L_0_out : std_logic := '0'; 
signal C_10_S_1_L_1_out : std_logic := '0'; 
signal C_10_S_1_L_2_out : std_logic := '0'; 
signal C_10_S_1_L_3_out : std_logic := '0'; 
signal C_10_S_1_L_4_out : std_logic := '0'; 
signal C_10_S_1_L_5_out : std_logic := '0'; 
signal C_10_S_2_L_0_out : std_logic := '0'; 
signal C_10_S_2_L_1_out : std_logic := '0'; 
signal C_10_S_2_L_2_out : std_logic := '0'; 
signal C_10_S_2_L_3_out : std_logic := '0'; 
signal C_10_S_2_L_4_out : std_logic := '0'; 
signal C_10_S_2_L_5_out : std_logic := '0'; 
signal C_10_S_3_L_0_out : std_logic := '0'; 
signal C_10_S_3_L_1_out : std_logic := '0'; 
signal C_10_S_3_L_2_out : std_logic := '0'; 
signal C_10_S_3_L_3_out : std_logic := '0'; 
signal C_10_S_3_L_4_out : std_logic := '0'; 
signal C_10_S_3_L_5_out : std_logic := '0'; 
signal C_10_S_4_L_0_out : std_logic := '0'; 
signal C_10_S_4_L_1_out : std_logic := '0'; 
signal C_10_S_4_L_2_out : std_logic := '0'; 
signal C_10_S_4_L_3_out : std_logic := '0'; 
signal C_10_S_4_L_4_out : std_logic := '0'; 
signal C_10_S_4_L_5_out : std_logic := '0'; 
signal C_10_S_5_L_0_out : std_logic := '0'; 
signal C_10_S_5_L_1_out : std_logic := '0'; 
signal C_10_S_5_L_2_out : std_logic := '0'; 
signal C_10_S_5_L_3_out : std_logic := '0'; 
signal C_10_S_5_L_4_out : std_logic := '0'; 
signal C_10_S_5_L_5_out : std_logic := '0'; 
signal C_11_S_0_L_0_out : std_logic := '0'; 
signal C_11_S_0_L_1_out : std_logic := '0'; 
signal C_11_S_0_L_2_out : std_logic := '0'; 
signal C_11_S_0_L_3_out : std_logic := '0'; 
signal C_11_S_0_L_4_out : std_logic := '0'; 
signal C_11_S_0_L_5_out : std_logic := '0'; 
signal C_11_S_1_L_0_out : std_logic := '0'; 
signal C_11_S_1_L_1_out : std_logic := '0'; 
signal C_11_S_1_L_2_out : std_logic := '0'; 
signal C_11_S_1_L_3_out : std_logic := '0'; 
signal C_11_S_1_L_4_out : std_logic := '0'; 
signal C_11_S_1_L_5_out : std_logic := '0'; 
signal C_11_S_2_L_0_out : std_logic := '0'; 
signal C_11_S_2_L_1_out : std_logic := '0'; 
signal C_11_S_2_L_2_out : std_logic := '0'; 
signal C_11_S_2_L_3_out : std_logic := '0'; 
signal C_11_S_2_L_4_out : std_logic := '0'; 
signal C_11_S_2_L_5_out : std_logic := '0'; 
signal C_11_S_3_L_0_out : std_logic := '0'; 
signal C_11_S_3_L_1_out : std_logic := '0'; 
signal C_11_S_3_L_2_out : std_logic := '0'; 
signal C_11_S_3_L_3_out : std_logic := '0'; 
signal C_11_S_3_L_4_out : std_logic := '0'; 
signal C_11_S_3_L_5_out : std_logic := '0'; 
signal C_11_S_4_L_0_out : std_logic := '0'; 
signal C_11_S_4_L_1_out : std_logic := '0'; 
signal C_11_S_4_L_2_out : std_logic := '0'; 
signal C_11_S_4_L_3_out : std_logic := '0'; 
signal C_11_S_4_L_4_out : std_logic := '0'; 
signal C_11_S_4_L_5_out : std_logic := '0'; 
signal C_11_S_5_L_0_out : std_logic := '0'; 
signal C_11_S_5_L_1_out : std_logic := '0'; 
signal C_11_S_5_L_2_out : std_logic := '0'; 
signal C_11_S_5_L_3_out : std_logic := '0'; 
signal C_11_S_5_L_4_out : std_logic := '0'; 
signal C_11_S_5_L_5_out : std_logic := '0'; 
signal C_12_S_0_L_0_out : std_logic := '0'; 
signal C_12_S_0_L_1_out : std_logic := '0'; 
signal C_12_S_0_L_2_out : std_logic := '0'; 
signal C_12_S_0_L_3_out : std_logic := '0'; 
signal C_12_S_0_L_4_out : std_logic := '0'; 
signal C_12_S_0_L_5_out : std_logic := '0'; 
signal C_12_S_1_L_0_out : std_logic := '0'; 
signal C_12_S_1_L_1_out : std_logic := '0'; 
signal C_12_S_1_L_2_out : std_logic := '0'; 
signal C_12_S_1_L_3_out : std_logic := '0'; 
signal C_12_S_1_L_4_out : std_logic := '0'; 
signal C_12_S_1_L_5_out : std_logic := '0'; 
signal C_12_S_2_L_0_out : std_logic := '0'; 
signal C_12_S_2_L_1_out : std_logic := '0'; 
signal C_12_S_2_L_2_out : std_logic := '0'; 
signal C_12_S_2_L_3_out : std_logic := '0'; 
signal C_12_S_2_L_4_out : std_logic := '0'; 
signal C_12_S_2_L_5_out : std_logic := '0'; 
signal C_12_S_3_L_0_out : std_logic := '0'; 
signal C_12_S_3_L_1_out : std_logic := '0'; 
signal C_12_S_3_L_2_out : std_logic := '0'; 
signal C_12_S_3_L_3_out : std_logic := '0'; 
signal C_12_S_3_L_4_out : std_logic := '0'; 
signal C_12_S_3_L_5_out : std_logic := '0'; 
signal C_12_S_4_L_0_out : std_logic := '0'; 
signal C_12_S_4_L_1_out : std_logic := '0'; 
signal C_12_S_4_L_2_out : std_logic := '0'; 
signal C_12_S_4_L_3_out : std_logic := '0'; 
signal C_12_S_4_L_4_out : std_logic := '0'; 
signal C_12_S_4_L_5_out : std_logic := '0'; 
signal C_12_S_5_L_0_out : std_logic := '0'; 
signal C_12_S_5_L_1_out : std_logic := '0'; 
signal C_12_S_5_L_2_out : std_logic := '0'; 
signal C_12_S_5_L_3_out : std_logic := '0'; 
signal C_12_S_5_L_4_out : std_logic := '0'; 
signal C_12_S_5_L_5_out : std_logic := '0'; 
signal C_13_S_0_L_0_out : std_logic := '0'; 
signal C_13_S_0_L_1_out : std_logic := '0'; 
signal C_13_S_0_L_2_out : std_logic := '0'; 
signal C_13_S_0_L_3_out : std_logic := '0'; 
signal C_13_S_0_L_4_out : std_logic := '0'; 
signal C_13_S_0_L_5_out : std_logic := '0'; 
signal C_13_S_1_L_0_out : std_logic := '0'; 
signal C_13_S_1_L_1_out : std_logic := '0'; 
signal C_13_S_1_L_2_out : std_logic := '0'; 
signal C_13_S_1_L_3_out : std_logic := '0'; 
signal C_13_S_1_L_4_out : std_logic := '0'; 
signal C_13_S_1_L_5_out : std_logic := '0'; 
signal C_13_S_2_L_0_out : std_logic := '0'; 
signal C_13_S_2_L_1_out : std_logic := '0'; 
signal C_13_S_2_L_2_out : std_logic := '0'; 
signal C_13_S_2_L_3_out : std_logic := '0'; 
signal C_13_S_2_L_4_out : std_logic := '0'; 
signal C_13_S_2_L_5_out : std_logic := '0'; 
signal C_13_S_3_L_0_out : std_logic := '0'; 
signal C_13_S_3_L_1_out : std_logic := '0'; 
signal C_13_S_3_L_2_out : std_logic := '0'; 
signal C_13_S_3_L_3_out : std_logic := '0'; 
signal C_13_S_3_L_4_out : std_logic := '0'; 
signal C_13_S_3_L_5_out : std_logic := '0'; 
signal C_13_S_4_L_0_out : std_logic := '0'; 
signal C_13_S_4_L_1_out : std_logic := '0'; 
signal C_13_S_4_L_2_out : std_logic := '0'; 
signal C_13_S_4_L_3_out : std_logic := '0'; 
signal C_13_S_4_L_4_out : std_logic := '0'; 
signal C_13_S_4_L_5_out : std_logic := '0'; 
signal C_13_S_5_L_0_out : std_logic := '0'; 
signal C_13_S_5_L_1_out : std_logic := '0'; 
signal C_13_S_5_L_2_out : std_logic := '0'; 
signal C_13_S_5_L_3_out : std_logic := '0'; 
signal C_13_S_5_L_4_out : std_logic := '0'; 
signal C_13_S_5_L_5_out : std_logic := '0'; 
signal C_14_S_0_L_0_out : std_logic := '0'; 
signal C_14_S_0_L_1_out : std_logic := '0'; 
signal C_14_S_0_L_2_out : std_logic := '0'; 
signal C_14_S_0_L_3_out : std_logic := '0'; 
signal C_14_S_0_L_4_out : std_logic := '0'; 
signal C_14_S_0_L_5_out : std_logic := '0'; 
signal C_14_S_1_L_0_out : std_logic := '0'; 
signal C_14_S_1_L_1_out : std_logic := '0'; 
signal C_14_S_1_L_2_out : std_logic := '0'; 
signal C_14_S_1_L_3_out : std_logic := '0'; 
signal C_14_S_1_L_4_out : std_logic := '0'; 
signal C_14_S_1_L_5_out : std_logic := '0'; 
signal C_14_S_2_L_0_out : std_logic := '0'; 
signal C_14_S_2_L_1_out : std_logic := '0'; 
signal C_14_S_2_L_2_out : std_logic := '0'; 
signal C_14_S_2_L_3_out : std_logic := '0'; 
signal C_14_S_2_L_4_out : std_logic := '0'; 
signal C_14_S_2_L_5_out : std_logic := '0'; 
signal C_14_S_3_L_0_out : std_logic := '0'; 
signal C_14_S_3_L_1_out : std_logic := '0'; 
signal C_14_S_3_L_2_out : std_logic := '0'; 
signal C_14_S_3_L_3_out : std_logic := '0'; 
signal C_14_S_3_L_4_out : std_logic := '0'; 
signal C_14_S_3_L_5_out : std_logic := '0'; 
signal C_14_S_4_L_0_out : std_logic := '0'; 
signal C_14_S_4_L_1_out : std_logic := '0'; 
signal C_14_S_4_L_2_out : std_logic := '0'; 
signal C_14_S_4_L_3_out : std_logic := '0'; 
signal C_14_S_4_L_4_out : std_logic := '0'; 
signal C_14_S_4_L_5_out : std_logic := '0'; 
signal C_14_S_5_L_0_out : std_logic := '0'; 
signal C_14_S_5_L_1_out : std_logic := '0'; 
signal C_14_S_5_L_2_out : std_logic := '0'; 
signal C_14_S_5_L_3_out : std_logic := '0'; 
signal C_14_S_5_L_4_out : std_logic := '0'; 
signal C_14_S_5_L_5_out : std_logic := '0'; 
signal C_15_S_0_L_0_out : std_logic := '0'; 
signal C_15_S_0_L_1_out : std_logic := '0'; 
signal C_15_S_0_L_2_out : std_logic := '0'; 
signal C_15_S_0_L_3_out : std_logic := '0'; 
signal C_15_S_0_L_4_out : std_logic := '0'; 
signal C_15_S_0_L_5_out : std_logic := '0'; 
signal C_15_S_1_L_0_out : std_logic := '0'; 
signal C_15_S_1_L_1_out : std_logic := '0'; 
signal C_15_S_1_L_2_out : std_logic := '0'; 
signal C_15_S_1_L_3_out : std_logic := '0'; 
signal C_15_S_1_L_4_out : std_logic := '0'; 
signal C_15_S_1_L_5_out : std_logic := '0'; 
signal C_15_S_2_L_0_out : std_logic := '0'; 
signal C_15_S_2_L_1_out : std_logic := '0'; 
signal C_15_S_2_L_2_out : std_logic := '0'; 
signal C_15_S_2_L_3_out : std_logic := '0'; 
signal C_15_S_2_L_4_out : std_logic := '0'; 
signal C_15_S_2_L_5_out : std_logic := '0'; 
signal C_15_S_3_L_0_out : std_logic := '0'; 
signal C_15_S_3_L_1_out : std_logic := '0'; 
signal C_15_S_3_L_2_out : std_logic := '0'; 
signal C_15_S_3_L_3_out : std_logic := '0'; 
signal C_15_S_3_L_4_out : std_logic := '0'; 
signal C_15_S_3_L_5_out : std_logic := '0'; 
signal C_15_S_4_L_0_out : std_logic := '0'; 
signal C_15_S_4_L_1_out : std_logic := '0'; 
signal C_15_S_4_L_2_out : std_logic := '0'; 
signal C_15_S_4_L_3_out : std_logic := '0'; 
signal C_15_S_4_L_4_out : std_logic := '0'; 
signal C_15_S_4_L_5_out : std_logic := '0'; 
signal C_15_S_5_L_0_out : std_logic := '0'; 
signal C_15_S_5_L_1_out : std_logic := '0'; 
signal C_15_S_5_L_2_out : std_logic := '0'; 
signal C_15_S_5_L_3_out : std_logic := '0'; 
signal C_15_S_5_L_4_out : std_logic := '0'; 
signal C_15_S_5_L_5_out : std_logic := '0'; 
signal C_16_S_0_L_0_out : std_logic := '0'; 
signal C_16_S_0_L_1_out : std_logic := '0'; 
signal C_16_S_0_L_2_out : std_logic := '0'; 
signal C_16_S_0_L_3_out : std_logic := '0'; 
signal C_16_S_0_L_4_out : std_logic := '0'; 
signal C_16_S_0_L_5_out : std_logic := '0'; 
signal C_16_S_1_L_0_out : std_logic := '0'; 
signal C_16_S_1_L_1_out : std_logic := '0'; 
signal C_16_S_1_L_2_out : std_logic := '0'; 
signal C_16_S_1_L_3_out : std_logic := '0'; 
signal C_16_S_1_L_4_out : std_logic := '0'; 
signal C_16_S_1_L_5_out : std_logic := '0'; 
signal C_16_S_2_L_0_out : std_logic := '0'; 
signal C_16_S_2_L_1_out : std_logic := '0'; 
signal C_16_S_2_L_2_out : std_logic := '0'; 
signal C_16_S_2_L_3_out : std_logic := '0'; 
signal C_16_S_2_L_4_out : std_logic := '0'; 
signal C_16_S_2_L_5_out : std_logic := '0'; 
signal C_16_S_3_L_0_out : std_logic := '0'; 
signal C_16_S_3_L_1_out : std_logic := '0'; 
signal C_16_S_3_L_2_out : std_logic := '0'; 
signal C_16_S_3_L_3_out : std_logic := '0'; 
signal C_16_S_3_L_4_out : std_logic := '0'; 
signal C_16_S_3_L_5_out : std_logic := '0'; 
signal C_16_S_4_L_0_out : std_logic := '0'; 
signal C_16_S_4_L_1_out : std_logic := '0'; 
signal C_16_S_4_L_2_out : std_logic := '0'; 
signal C_16_S_4_L_3_out : std_logic := '0'; 
signal C_16_S_4_L_4_out : std_logic := '0'; 
signal C_16_S_4_L_5_out : std_logic := '0'; 
signal C_16_S_5_L_0_out : std_logic := '0'; 
signal C_16_S_5_L_1_out : std_logic := '0'; 
signal C_16_S_5_L_2_out : std_logic := '0'; 
signal C_16_S_5_L_3_out : std_logic := '0'; 
signal C_16_S_5_L_4_out : std_logic := '0'; 
signal C_16_S_5_L_5_out : std_logic := '0'; 
signal C_17_S_0_L_0_out : std_logic := '0'; 
signal C_17_S_0_L_1_out : std_logic := '0'; 
signal C_17_S_0_L_2_out : std_logic := '0'; 
signal C_17_S_0_L_3_out : std_logic := '0'; 
signal C_17_S_0_L_4_out : std_logic := '0'; 
signal C_17_S_0_L_5_out : std_logic := '0'; 
signal C_17_S_1_L_0_out : std_logic := '0'; 
signal C_17_S_1_L_1_out : std_logic := '0'; 
signal C_17_S_1_L_2_out : std_logic := '0'; 
signal C_17_S_1_L_3_out : std_logic := '0'; 
signal C_17_S_1_L_4_out : std_logic := '0'; 
signal C_17_S_1_L_5_out : std_logic := '0'; 
signal C_17_S_2_L_0_out : std_logic := '0'; 
signal C_17_S_2_L_1_out : std_logic := '0'; 
signal C_17_S_2_L_2_out : std_logic := '0'; 
signal C_17_S_2_L_3_out : std_logic := '0'; 
signal C_17_S_2_L_4_out : std_logic := '0'; 
signal C_17_S_2_L_5_out : std_logic := '0'; 
signal C_17_S_3_L_0_out : std_logic := '0'; 
signal C_17_S_3_L_1_out : std_logic := '0'; 
signal C_17_S_3_L_2_out : std_logic := '0'; 
signal C_17_S_3_L_3_out : std_logic := '0'; 
signal C_17_S_3_L_4_out : std_logic := '0'; 
signal C_17_S_3_L_5_out : std_logic := '0'; 
signal C_17_S_4_L_0_out : std_logic := '0'; 
signal C_17_S_4_L_1_out : std_logic := '0'; 
signal C_17_S_4_L_2_out : std_logic := '0'; 
signal C_17_S_4_L_3_out : std_logic := '0'; 
signal C_17_S_4_L_4_out : std_logic := '0'; 
signal C_17_S_4_L_5_out : std_logic := '0'; 
signal C_17_S_5_L_0_out : std_logic := '0'; 
signal C_17_S_5_L_1_out : std_logic := '0'; 
signal C_17_S_5_L_2_out : std_logic := '0'; 
signal C_17_S_5_L_3_out : std_logic := '0'; 
signal C_17_S_5_L_4_out : std_logic := '0'; 
signal C_17_S_5_L_5_out : std_logic := '0'; 
signal C_18_S_0_L_0_out : std_logic := '0'; 
signal C_18_S_0_L_1_out : std_logic := '0'; 
signal C_18_S_0_L_2_out : std_logic := '0'; 
signal C_18_S_0_L_3_out : std_logic := '0'; 
signal C_18_S_0_L_4_out : std_logic := '0'; 
signal C_18_S_0_L_5_out : std_logic := '0'; 
signal C_18_S_1_L_0_out : std_logic := '0'; 
signal C_18_S_1_L_1_out : std_logic := '0'; 
signal C_18_S_1_L_2_out : std_logic := '0'; 
signal C_18_S_1_L_3_out : std_logic := '0'; 
signal C_18_S_1_L_4_out : std_logic := '0'; 
signal C_18_S_1_L_5_out : std_logic := '0'; 
signal C_18_S_2_L_0_out : std_logic := '0'; 
signal C_18_S_2_L_1_out : std_logic := '0'; 
signal C_18_S_2_L_2_out : std_logic := '0'; 
signal C_18_S_2_L_3_out : std_logic := '0'; 
signal C_18_S_2_L_4_out : std_logic := '0'; 
signal C_18_S_2_L_5_out : std_logic := '0'; 
signal C_18_S_3_L_0_out : std_logic := '0'; 
signal C_18_S_3_L_1_out : std_logic := '0'; 
signal C_18_S_3_L_2_out : std_logic := '0'; 
signal C_18_S_3_L_3_out : std_logic := '0'; 
signal C_18_S_3_L_4_out : std_logic := '0'; 
signal C_18_S_3_L_5_out : std_logic := '0'; 
signal C_18_S_4_L_0_out : std_logic := '0'; 
signal C_18_S_4_L_1_out : std_logic := '0'; 
signal C_18_S_4_L_2_out : std_logic := '0'; 
signal C_18_S_4_L_3_out : std_logic := '0'; 
signal C_18_S_4_L_4_out : std_logic := '0'; 
signal C_18_S_4_L_5_out : std_logic := '0'; 
signal C_18_S_5_L_0_out : std_logic := '0'; 
signal C_18_S_5_L_1_out : std_logic := '0'; 
signal C_18_S_5_L_2_out : std_logic := '0'; 
signal C_18_S_5_L_3_out : std_logic := '0'; 
signal C_18_S_5_L_4_out : std_logic := '0'; 
signal C_18_S_5_L_5_out : std_logic := '0'; 
signal C_19_S_0_L_0_out : std_logic := '0'; 
signal C_19_S_0_L_1_out : std_logic := '0'; 
signal C_19_S_0_L_2_out : std_logic := '0'; 
signal C_19_S_0_L_3_out : std_logic := '0'; 
signal C_19_S_0_L_4_out : std_logic := '0'; 
signal C_19_S_0_L_5_out : std_logic := '0'; 
signal C_19_S_1_L_0_out : std_logic := '0'; 
signal C_19_S_1_L_1_out : std_logic := '0'; 
signal C_19_S_1_L_2_out : std_logic := '0'; 
signal C_19_S_1_L_3_out : std_logic := '0'; 
signal C_19_S_1_L_4_out : std_logic := '0'; 
signal C_19_S_1_L_5_out : std_logic := '0'; 
signal C_19_S_2_L_0_out : std_logic := '0'; 
signal C_19_S_2_L_1_out : std_logic := '0'; 
signal C_19_S_2_L_2_out : std_logic := '0'; 
signal C_19_S_2_L_3_out : std_logic := '0'; 
signal C_19_S_2_L_4_out : std_logic := '0'; 
signal C_19_S_2_L_5_out : std_logic := '0'; 
signal C_19_S_3_L_0_out : std_logic := '0'; 
signal C_19_S_3_L_1_out : std_logic := '0'; 
signal C_19_S_3_L_2_out : std_logic := '0'; 
signal C_19_S_3_L_3_out : std_logic := '0'; 
signal C_19_S_3_L_4_out : std_logic := '0'; 
signal C_19_S_3_L_5_out : std_logic := '0'; 
signal C_19_S_4_L_0_out : std_logic := '0'; 
signal C_19_S_4_L_1_out : std_logic := '0'; 
signal C_19_S_4_L_2_out : std_logic := '0'; 
signal C_19_S_4_L_3_out : std_logic := '0'; 
signal C_19_S_4_L_4_out : std_logic := '0'; 
signal C_19_S_4_L_5_out : std_logic := '0'; 
signal C_19_S_5_L_0_out : std_logic := '0'; 
signal C_19_S_5_L_1_out : std_logic := '0'; 
signal C_19_S_5_L_2_out : std_logic := '0'; 
signal C_19_S_5_L_3_out : std_logic := '0'; 
signal C_19_S_5_L_4_out : std_logic := '0'; 
signal C_19_S_5_L_5_out : std_logic := '0'; 
signal C_20_S_0_L_0_out : std_logic := '0'; 
signal C_20_S_0_L_1_out : std_logic := '0'; 
signal C_20_S_0_L_2_out : std_logic := '0'; 
signal C_20_S_0_L_3_out : std_logic := '0'; 
signal C_20_S_0_L_4_out : std_logic := '0'; 
signal C_20_S_0_L_5_out : std_logic := '0'; 
signal C_20_S_1_L_0_out : std_logic := '0'; 
signal C_20_S_1_L_1_out : std_logic := '0'; 
signal C_20_S_1_L_2_out : std_logic := '0'; 
signal C_20_S_1_L_3_out : std_logic := '0'; 
signal C_20_S_1_L_4_out : std_logic := '0'; 
signal C_20_S_1_L_5_out : std_logic := '0'; 
signal C_20_S_2_L_0_out : std_logic := '0'; 
signal C_20_S_2_L_1_out : std_logic := '0'; 
signal C_20_S_2_L_2_out : std_logic := '0'; 
signal C_20_S_2_L_3_out : std_logic := '0'; 
signal C_20_S_2_L_4_out : std_logic := '0'; 
signal C_20_S_2_L_5_out : std_logic := '0'; 
signal C_20_S_3_L_0_out : std_logic := '0'; 
signal C_20_S_3_L_1_out : std_logic := '0'; 
signal C_20_S_3_L_2_out : std_logic := '0'; 
signal C_20_S_3_L_3_out : std_logic := '0'; 
signal C_20_S_3_L_4_out : std_logic := '0'; 
signal C_20_S_3_L_5_out : std_logic := '0'; 
signal C_20_S_4_L_0_out : std_logic := '0'; 
signal C_20_S_4_L_1_out : std_logic := '0'; 
signal C_20_S_4_L_2_out : std_logic := '0'; 
signal C_20_S_4_L_3_out : std_logic := '0'; 
signal C_20_S_4_L_4_out : std_logic := '0'; 
signal C_20_S_4_L_5_out : std_logic := '0'; 
signal C_20_S_5_L_0_out : std_logic := '0'; 
signal C_20_S_5_L_1_out : std_logic := '0'; 
signal C_20_S_5_L_2_out : std_logic := '0'; 
signal C_20_S_5_L_3_out : std_logic := '0'; 
signal C_20_S_5_L_4_out : std_logic := '0'; 
signal C_20_S_5_L_5_out : std_logic := '0'; 
signal C_21_S_0_L_0_out : std_logic := '0'; 
signal C_21_S_0_L_1_out : std_logic := '0'; 
signal C_21_S_0_L_2_out : std_logic := '0'; 
signal C_21_S_0_L_3_out : std_logic := '0'; 
signal C_21_S_0_L_4_out : std_logic := '0'; 
signal C_21_S_0_L_5_out : std_logic := '0'; 
signal C_21_S_1_L_0_out : std_logic := '0'; 
signal C_21_S_1_L_1_out : std_logic := '0'; 
signal C_21_S_1_L_2_out : std_logic := '0'; 
signal C_21_S_1_L_3_out : std_logic := '0'; 
signal C_21_S_1_L_4_out : std_logic := '0'; 
signal C_21_S_1_L_5_out : std_logic := '0'; 
signal C_21_S_2_L_0_out : std_logic := '0'; 
signal C_21_S_2_L_1_out : std_logic := '0'; 
signal C_21_S_2_L_2_out : std_logic := '0'; 
signal C_21_S_2_L_3_out : std_logic := '0'; 
signal C_21_S_2_L_4_out : std_logic := '0'; 
signal C_21_S_2_L_5_out : std_logic := '0'; 
signal C_21_S_3_L_0_out : std_logic := '0'; 
signal C_21_S_3_L_1_out : std_logic := '0'; 
signal C_21_S_3_L_2_out : std_logic := '0'; 
signal C_21_S_3_L_3_out : std_logic := '0'; 
signal C_21_S_3_L_4_out : std_logic := '0'; 
signal C_21_S_3_L_5_out : std_logic := '0'; 
signal C_21_S_4_L_0_out : std_logic := '0'; 
signal C_21_S_4_L_1_out : std_logic := '0'; 
signal C_21_S_4_L_2_out : std_logic := '0'; 
signal C_21_S_4_L_3_out : std_logic := '0'; 
signal C_21_S_4_L_4_out : std_logic := '0'; 
signal C_21_S_4_L_5_out : std_logic := '0'; 
signal C_21_S_5_L_0_out : std_logic := '0'; 
signal C_21_S_5_L_1_out : std_logic := '0'; 
signal C_21_S_5_L_2_out : std_logic := '0'; 
signal C_21_S_5_L_3_out : std_logic := '0'; 
signal C_21_S_5_L_4_out : std_logic := '0'; 
signal C_21_S_5_L_5_out : std_logic := '0'; 
signal C_22_S_0_L_0_out : std_logic := '0'; 
signal C_22_S_0_L_1_out : std_logic := '0'; 
signal C_22_S_0_L_2_out : std_logic := '0'; 
signal C_22_S_0_L_3_out : std_logic := '0'; 
signal C_22_S_0_L_4_out : std_logic := '0'; 
signal C_22_S_0_L_5_out : std_logic := '0'; 
signal C_22_S_1_L_0_out : std_logic := '0'; 
signal C_22_S_1_L_1_out : std_logic := '0'; 
signal C_22_S_1_L_2_out : std_logic := '0'; 
signal C_22_S_1_L_3_out : std_logic := '0'; 
signal C_22_S_1_L_4_out : std_logic := '0'; 
signal C_22_S_1_L_5_out : std_logic := '0'; 
signal C_22_S_2_L_0_out : std_logic := '0'; 
signal C_22_S_2_L_1_out : std_logic := '0'; 
signal C_22_S_2_L_2_out : std_logic := '0'; 
signal C_22_S_2_L_3_out : std_logic := '0'; 
signal C_22_S_2_L_4_out : std_logic := '0'; 
signal C_22_S_2_L_5_out : std_logic := '0'; 
signal C_22_S_3_L_0_out : std_logic := '0'; 
signal C_22_S_3_L_1_out : std_logic := '0'; 
signal C_22_S_3_L_2_out : std_logic := '0'; 
signal C_22_S_3_L_3_out : std_logic := '0'; 
signal C_22_S_3_L_4_out : std_logic := '0'; 
signal C_22_S_3_L_5_out : std_logic := '0'; 
signal C_22_S_4_L_0_out : std_logic := '0'; 
signal C_22_S_4_L_1_out : std_logic := '0'; 
signal C_22_S_4_L_2_out : std_logic := '0'; 
signal C_22_S_4_L_3_out : std_logic := '0'; 
signal C_22_S_4_L_4_out : std_logic := '0'; 
signal C_22_S_4_L_5_out : std_logic := '0'; 
signal C_22_S_5_L_0_out : std_logic := '0'; 
signal C_22_S_5_L_1_out : std_logic := '0'; 
signal C_22_S_5_L_2_out : std_logic := '0'; 
signal C_22_S_5_L_3_out : std_logic := '0'; 
signal C_22_S_5_L_4_out : std_logic := '0'; 
signal C_22_S_5_L_5_out : std_logic := '0'; 
signal C_23_S_0_L_0_out : std_logic := '0'; 
signal C_23_S_0_L_1_out : std_logic := '0'; 
signal C_23_S_0_L_2_out : std_logic := '0'; 
signal C_23_S_0_L_3_out : std_logic := '0'; 
signal C_23_S_0_L_4_out : std_logic := '0'; 
signal C_23_S_0_L_5_out : std_logic := '0'; 
signal C_23_S_1_L_0_out : std_logic := '0'; 
signal C_23_S_1_L_1_out : std_logic := '0'; 
signal C_23_S_1_L_2_out : std_logic := '0'; 
signal C_23_S_1_L_3_out : std_logic := '0'; 
signal C_23_S_1_L_4_out : std_logic := '0'; 
signal C_23_S_1_L_5_out : std_logic := '0'; 
signal C_23_S_2_L_0_out : std_logic := '0'; 
signal C_23_S_2_L_1_out : std_logic := '0'; 
signal C_23_S_2_L_2_out : std_logic := '0'; 
signal C_23_S_2_L_3_out : std_logic := '0'; 
signal C_23_S_2_L_4_out : std_logic := '0'; 
signal C_23_S_2_L_5_out : std_logic := '0'; 
signal C_23_S_3_L_0_out : std_logic := '0'; 
signal C_23_S_3_L_1_out : std_logic := '0'; 
signal C_23_S_3_L_2_out : std_logic := '0'; 
signal C_23_S_3_L_3_out : std_logic := '0'; 
signal C_23_S_3_L_4_out : std_logic := '0'; 
signal C_23_S_3_L_5_out : std_logic := '0'; 
signal C_23_S_4_L_0_out : std_logic := '0'; 
signal C_23_S_4_L_1_out : std_logic := '0'; 
signal C_23_S_4_L_2_out : std_logic := '0'; 
signal C_23_S_4_L_3_out : std_logic := '0'; 
signal C_23_S_4_L_4_out : std_logic := '0'; 
signal C_23_S_4_L_5_out : std_logic := '0'; 
signal C_23_S_5_L_0_out : std_logic := '0'; 
signal C_23_S_5_L_1_out : std_logic := '0'; 
signal C_23_S_5_L_2_out : std_logic := '0'; 
signal C_23_S_5_L_3_out : std_logic := '0'; 
signal C_23_S_5_L_4_out : std_logic := '0'; 
signal C_23_S_5_L_5_out : std_logic := '0'; 
signal C_24_S_0_L_0_out : std_logic := '0'; 
signal C_24_S_0_L_1_out : std_logic := '0'; 
signal C_24_S_0_L_2_out : std_logic := '0'; 
signal C_24_S_0_L_3_out : std_logic := '0'; 
signal C_24_S_0_L_4_out : std_logic := '0'; 
signal C_24_S_0_L_5_out : std_logic := '0'; 
signal C_24_S_1_L_0_out : std_logic := '0'; 
signal C_24_S_1_L_1_out : std_logic := '0'; 
signal C_24_S_1_L_2_out : std_logic := '0'; 
signal C_24_S_1_L_3_out : std_logic := '0'; 
signal C_24_S_1_L_4_out : std_logic := '0'; 
signal C_24_S_1_L_5_out : std_logic := '0'; 
signal C_24_S_2_L_0_out : std_logic := '0'; 
signal C_24_S_2_L_1_out : std_logic := '0'; 
signal C_24_S_2_L_2_out : std_logic := '0'; 
signal C_24_S_2_L_3_out : std_logic := '0'; 
signal C_24_S_2_L_4_out : std_logic := '0'; 
signal C_24_S_2_L_5_out : std_logic := '0'; 
signal C_24_S_3_L_0_out : std_logic := '0'; 
signal C_24_S_3_L_1_out : std_logic := '0'; 
signal C_24_S_3_L_2_out : std_logic := '0'; 
signal C_24_S_3_L_3_out : std_logic := '0'; 
signal C_24_S_3_L_4_out : std_logic := '0'; 
signal C_24_S_3_L_5_out : std_logic := '0'; 
signal C_24_S_4_L_0_out : std_logic := '0'; 
signal C_24_S_4_L_1_out : std_logic := '0'; 
signal C_24_S_4_L_2_out : std_logic := '0'; 
signal C_24_S_4_L_3_out : std_logic := '0'; 
signal C_24_S_4_L_4_out : std_logic := '0'; 
signal C_24_S_4_L_5_out : std_logic := '0'; 
signal C_24_S_5_L_0_out : std_logic := '0'; 
signal C_24_S_5_L_1_out : std_logic := '0'; 
signal C_24_S_5_L_2_out : std_logic := '0'; 
signal C_24_S_5_L_3_out : std_logic := '0'; 
signal C_24_S_5_L_4_out : std_logic := '0'; 
signal C_24_S_5_L_5_out : std_logic := '0'; 
signal C_25_S_0_L_0_out : std_logic := '0'; 
signal C_25_S_0_L_1_out : std_logic := '0'; 
signal C_25_S_0_L_2_out : std_logic := '0'; 
signal C_25_S_0_L_3_out : std_logic := '0'; 
signal C_25_S_0_L_4_out : std_logic := '0'; 
signal C_25_S_0_L_5_out : std_logic := '0'; 
signal C_25_S_1_L_0_out : std_logic := '0'; 
signal C_25_S_1_L_1_out : std_logic := '0'; 
signal C_25_S_1_L_2_out : std_logic := '0'; 
signal C_25_S_1_L_3_out : std_logic := '0'; 
signal C_25_S_1_L_4_out : std_logic := '0'; 
signal C_25_S_1_L_5_out : std_logic := '0'; 
signal C_25_S_2_L_0_out : std_logic := '0'; 
signal C_25_S_2_L_1_out : std_logic := '0'; 
signal C_25_S_2_L_2_out : std_logic := '0'; 
signal C_25_S_2_L_3_out : std_logic := '0'; 
signal C_25_S_2_L_4_out : std_logic := '0'; 
signal C_25_S_2_L_5_out : std_logic := '0'; 
signal C_25_S_3_L_0_out : std_logic := '0'; 
signal C_25_S_3_L_1_out : std_logic := '0'; 
signal C_25_S_3_L_2_out : std_logic := '0'; 
signal C_25_S_3_L_3_out : std_logic := '0'; 
signal C_25_S_3_L_4_out : std_logic := '0'; 
signal C_25_S_3_L_5_out : std_logic := '0'; 
signal C_25_S_4_L_0_out : std_logic := '0'; 
signal C_25_S_4_L_1_out : std_logic := '0'; 
signal C_25_S_4_L_2_out : std_logic := '0'; 
signal C_25_S_4_L_3_out : std_logic := '0'; 
signal C_25_S_4_L_4_out : std_logic := '0'; 
signal C_25_S_4_L_5_out : std_logic := '0'; 
signal C_25_S_5_L_0_out : std_logic := '0'; 
signal C_25_S_5_L_1_out : std_logic := '0'; 
signal C_25_S_5_L_2_out : std_logic := '0'; 
signal C_25_S_5_L_3_out : std_logic := '0'; 
signal C_25_S_5_L_4_out : std_logic := '0'; 
signal C_25_S_5_L_5_out : std_logic := '0'; 
signal C_26_S_0_L_0_out : std_logic := '0'; 
signal C_26_S_0_L_1_out : std_logic := '0'; 
signal C_26_S_0_L_2_out : std_logic := '0'; 
signal C_26_S_0_L_3_out : std_logic := '0'; 
signal C_26_S_0_L_4_out : std_logic := '0'; 
signal C_26_S_0_L_5_out : std_logic := '0'; 
signal C_26_S_1_L_0_out : std_logic := '0'; 
signal C_26_S_1_L_1_out : std_logic := '0'; 
signal C_26_S_1_L_2_out : std_logic := '0'; 
signal C_26_S_1_L_3_out : std_logic := '0'; 
signal C_26_S_1_L_4_out : std_logic := '0'; 
signal C_26_S_1_L_5_out : std_logic := '0'; 
signal C_26_S_2_L_0_out : std_logic := '0'; 
signal C_26_S_2_L_1_out : std_logic := '0'; 
signal C_26_S_2_L_2_out : std_logic := '0'; 
signal C_26_S_2_L_3_out : std_logic := '0'; 
signal C_26_S_2_L_4_out : std_logic := '0'; 
signal C_26_S_2_L_5_out : std_logic := '0'; 
signal C_26_S_3_L_0_out : std_logic := '0'; 
signal C_26_S_3_L_1_out : std_logic := '0'; 
signal C_26_S_3_L_2_out : std_logic := '0'; 
signal C_26_S_3_L_3_out : std_logic := '0'; 
signal C_26_S_3_L_4_out : std_logic := '0'; 
signal C_26_S_3_L_5_out : std_logic := '0'; 
signal C_26_S_4_L_0_out : std_logic := '0'; 
signal C_26_S_4_L_1_out : std_logic := '0'; 
signal C_26_S_4_L_2_out : std_logic := '0'; 
signal C_26_S_4_L_3_out : std_logic := '0'; 
signal C_26_S_4_L_4_out : std_logic := '0'; 
signal C_26_S_4_L_5_out : std_logic := '0'; 
signal C_26_S_5_L_0_out : std_logic := '0'; 
signal C_26_S_5_L_1_out : std_logic := '0'; 
signal C_26_S_5_L_2_out : std_logic := '0'; 
signal C_26_S_5_L_3_out : std_logic := '0'; 
signal C_26_S_5_L_4_out : std_logic := '0'; 
signal C_26_S_5_L_5_out : std_logic := '0'; 
signal C_27_S_0_L_0_out : std_logic := '0'; 
signal C_27_S_0_L_1_out : std_logic := '0'; 
signal C_27_S_0_L_2_out : std_logic := '0'; 
signal C_27_S_0_L_3_out : std_logic := '0'; 
signal C_27_S_0_L_4_out : std_logic := '0'; 
signal C_27_S_0_L_5_out : std_logic := '0'; 
signal C_27_S_1_L_0_out : std_logic := '0'; 
signal C_27_S_1_L_1_out : std_logic := '0'; 
signal C_27_S_1_L_2_out : std_logic := '0'; 
signal C_27_S_1_L_3_out : std_logic := '0'; 
signal C_27_S_1_L_4_out : std_logic := '0'; 
signal C_27_S_1_L_5_out : std_logic := '0'; 
signal C_27_S_2_L_0_out : std_logic := '0'; 
signal C_27_S_2_L_1_out : std_logic := '0'; 
signal C_27_S_2_L_2_out : std_logic := '0'; 
signal C_27_S_2_L_3_out : std_logic := '0'; 
signal C_27_S_2_L_4_out : std_logic := '0'; 
signal C_27_S_2_L_5_out : std_logic := '0'; 
signal C_27_S_3_L_0_out : std_logic := '0'; 
signal C_27_S_3_L_1_out : std_logic := '0'; 
signal C_27_S_3_L_2_out : std_logic := '0'; 
signal C_27_S_3_L_3_out : std_logic := '0'; 
signal C_27_S_3_L_4_out : std_logic := '0'; 
signal C_27_S_3_L_5_out : std_logic := '0'; 
signal C_27_S_4_L_0_out : std_logic := '0'; 
signal C_27_S_4_L_1_out : std_logic := '0'; 
signal C_27_S_4_L_2_out : std_logic := '0'; 
signal C_27_S_4_L_3_out : std_logic := '0'; 
signal C_27_S_4_L_4_out : std_logic := '0'; 
signal C_27_S_4_L_5_out : std_logic := '0'; 
signal C_27_S_5_L_0_out : std_logic := '0'; 
signal C_27_S_5_L_1_out : std_logic := '0'; 
signal C_27_S_5_L_2_out : std_logic := '0'; 
signal C_27_S_5_L_3_out : std_logic := '0'; 
signal C_27_S_5_L_4_out : std_logic := '0'; 
signal C_27_S_5_L_5_out : std_logic := '0'; 
signal C_28_S_0_L_0_out : std_logic := '0'; 
signal C_28_S_0_L_1_out : std_logic := '0'; 
signal C_28_S_0_L_2_out : std_logic := '0'; 
signal C_28_S_0_L_3_out : std_logic := '0'; 
signal C_28_S_0_L_4_out : std_logic := '0'; 
signal C_28_S_0_L_5_out : std_logic := '0'; 
signal C_28_S_1_L_0_out : std_logic := '0'; 
signal C_28_S_1_L_1_out : std_logic := '0'; 
signal C_28_S_1_L_2_out : std_logic := '0'; 
signal C_28_S_1_L_3_out : std_logic := '0'; 
signal C_28_S_1_L_4_out : std_logic := '0'; 
signal C_28_S_1_L_5_out : std_logic := '0'; 
signal C_28_S_2_L_0_out : std_logic := '0'; 
signal C_28_S_2_L_1_out : std_logic := '0'; 
signal C_28_S_2_L_2_out : std_logic := '0'; 
signal C_28_S_2_L_3_out : std_logic := '0'; 
signal C_28_S_2_L_4_out : std_logic := '0'; 
signal C_28_S_2_L_5_out : std_logic := '0'; 
signal C_28_S_3_L_0_out : std_logic := '0'; 
signal C_28_S_3_L_1_out : std_logic := '0'; 
signal C_28_S_3_L_2_out : std_logic := '0'; 
signal C_28_S_3_L_3_out : std_logic := '0'; 
signal C_28_S_3_L_4_out : std_logic := '0'; 
signal C_28_S_3_L_5_out : std_logic := '0'; 
signal C_28_S_4_L_0_out : std_logic := '0'; 
signal C_28_S_4_L_1_out : std_logic := '0'; 
signal C_28_S_4_L_2_out : std_logic := '0'; 
signal C_28_S_4_L_3_out : std_logic := '0'; 
signal C_28_S_4_L_4_out : std_logic := '0'; 
signal C_28_S_4_L_5_out : std_logic := '0'; 
signal C_28_S_5_L_0_out : std_logic := '0'; 
signal C_28_S_5_L_1_out : std_logic := '0'; 
signal C_28_S_5_L_2_out : std_logic := '0'; 
signal C_28_S_5_L_3_out : std_logic := '0'; 
signal C_28_S_5_L_4_out : std_logic := '0'; 
signal C_28_S_5_L_5_out : std_logic := '0'; 
signal C_29_S_0_L_0_out : std_logic := '0'; 
signal C_29_S_0_L_1_out : std_logic := '0'; 
signal C_29_S_0_L_2_out : std_logic := '0'; 
signal C_29_S_0_L_3_out : std_logic := '0'; 
signal C_29_S_0_L_4_out : std_logic := '0'; 
signal C_29_S_0_L_5_out : std_logic := '0'; 
signal C_29_S_1_L_0_out : std_logic := '0'; 
signal C_29_S_1_L_1_out : std_logic := '0'; 
signal C_29_S_1_L_2_out : std_logic := '0'; 
signal C_29_S_1_L_3_out : std_logic := '0'; 
signal C_29_S_1_L_4_out : std_logic := '0'; 
signal C_29_S_1_L_5_out : std_logic := '0'; 
signal C_29_S_2_L_0_out : std_logic := '0'; 
signal C_29_S_2_L_1_out : std_logic := '0'; 
signal C_29_S_2_L_2_out : std_logic := '0'; 
signal C_29_S_2_L_3_out : std_logic := '0'; 
signal C_29_S_2_L_4_out : std_logic := '0'; 
signal C_29_S_2_L_5_out : std_logic := '0'; 
signal C_29_S_3_L_0_out : std_logic := '0'; 
signal C_29_S_3_L_1_out : std_logic := '0'; 
signal C_29_S_3_L_2_out : std_logic := '0'; 
signal C_29_S_3_L_3_out : std_logic := '0'; 
signal C_29_S_3_L_4_out : std_logic := '0'; 
signal C_29_S_3_L_5_out : std_logic := '0'; 
signal C_29_S_4_L_0_out : std_logic := '0'; 
signal C_29_S_4_L_1_out : std_logic := '0'; 
signal C_29_S_4_L_2_out : std_logic := '0'; 
signal C_29_S_4_L_3_out : std_logic := '0'; 
signal C_29_S_4_L_4_out : std_logic := '0'; 
signal C_29_S_4_L_5_out : std_logic := '0'; 
signal C_29_S_5_L_0_out : std_logic := '0'; 
signal C_29_S_5_L_1_out : std_logic := '0'; 
signal C_29_S_5_L_2_out : std_logic := '0'; 
signal C_29_S_5_L_3_out : std_logic := '0'; 
signal C_29_S_5_L_4_out : std_logic := '0'; 
signal C_29_S_5_L_5_out : std_logic := '0'; 
signal C_30_S_0_L_0_out : std_logic := '0'; 
signal C_30_S_0_L_1_out : std_logic := '0'; 
signal C_30_S_0_L_2_out : std_logic := '0'; 
signal C_30_S_0_L_3_out : std_logic := '0'; 
signal C_30_S_0_L_4_out : std_logic := '0'; 
signal C_30_S_0_L_5_out : std_logic := '0'; 
signal C_30_S_1_L_0_out : std_logic := '0'; 
signal C_30_S_1_L_1_out : std_logic := '0'; 
signal C_30_S_1_L_2_out : std_logic := '0'; 
signal C_30_S_1_L_3_out : std_logic := '0'; 
signal C_30_S_1_L_4_out : std_logic := '0'; 
signal C_30_S_1_L_5_out : std_logic := '0'; 
signal C_30_S_2_L_0_out : std_logic := '0'; 
signal C_30_S_2_L_1_out : std_logic := '0'; 
signal C_30_S_2_L_2_out : std_logic := '0'; 
signal C_30_S_2_L_3_out : std_logic := '0'; 
signal C_30_S_2_L_4_out : std_logic := '0'; 
signal C_30_S_2_L_5_out : std_logic := '0'; 
signal C_30_S_3_L_0_out : std_logic := '0'; 
signal C_30_S_3_L_1_out : std_logic := '0'; 
signal C_30_S_3_L_2_out : std_logic := '0'; 
signal C_30_S_3_L_3_out : std_logic := '0'; 
signal C_30_S_3_L_4_out : std_logic := '0'; 
signal C_30_S_3_L_5_out : std_logic := '0'; 
signal C_30_S_4_L_0_out : std_logic := '0'; 
signal C_30_S_4_L_1_out : std_logic := '0'; 
signal C_30_S_4_L_2_out : std_logic := '0'; 
signal C_30_S_4_L_3_out : std_logic := '0'; 
signal C_30_S_4_L_4_out : std_logic := '0'; 
signal C_30_S_4_L_5_out : std_logic := '0'; 
signal C_30_S_5_L_0_out : std_logic := '0'; 
signal C_30_S_5_L_1_out : std_logic := '0'; 
signal C_30_S_5_L_2_out : std_logic := '0'; 
signal C_30_S_5_L_3_out : std_logic := '0'; 
signal C_30_S_5_L_4_out : std_logic := '0'; 
signal C_30_S_5_L_5_out : std_logic := '0'; 
signal C_31_S_0_L_0_out : std_logic := '0'; 
signal C_31_S_0_L_1_out : std_logic := '0'; 
signal C_31_S_0_L_2_out : std_logic := '0'; 
signal C_31_S_0_L_3_out : std_logic := '0'; 
signal C_31_S_0_L_4_out : std_logic := '0'; 
signal C_31_S_0_L_5_out : std_logic := '0'; 
signal C_31_S_1_L_0_out : std_logic := '0'; 
signal C_31_S_1_L_1_out : std_logic := '0'; 
signal C_31_S_1_L_2_out : std_logic := '0'; 
signal C_31_S_1_L_3_out : std_logic := '0'; 
signal C_31_S_1_L_4_out : std_logic := '0'; 
signal C_31_S_1_L_5_out : std_logic := '0'; 
signal C_31_S_2_L_0_out : std_logic := '0'; 
signal C_31_S_2_L_1_out : std_logic := '0'; 
signal C_31_S_2_L_2_out : std_logic := '0'; 
signal C_31_S_2_L_3_out : std_logic := '0'; 
signal C_31_S_2_L_4_out : std_logic := '0'; 
signal C_31_S_2_L_5_out : std_logic := '0'; 
signal C_31_S_3_L_0_out : std_logic := '0'; 
signal C_31_S_3_L_1_out : std_logic := '0'; 
signal C_31_S_3_L_2_out : std_logic := '0'; 
signal C_31_S_3_L_3_out : std_logic := '0'; 
signal C_31_S_3_L_4_out : std_logic := '0'; 
signal C_31_S_3_L_5_out : std_logic := '0'; 
signal C_31_S_4_L_0_out : std_logic := '0'; 
signal C_31_S_4_L_1_out : std_logic := '0'; 
signal C_31_S_4_L_2_out : std_logic := '0'; 
signal C_31_S_4_L_3_out : std_logic := '0'; 
signal C_31_S_4_L_4_out : std_logic := '0'; 
signal C_31_S_4_L_5_out : std_logic := '0'; 
signal C_31_S_5_L_0_out : std_logic := '0'; 
signal C_31_S_5_L_1_out : std_logic := '0'; 
signal C_31_S_5_L_2_out : std_logic := '0'; 
signal C_31_S_5_L_3_out : std_logic := '0'; 
signal C_31_S_5_L_4_out : std_logic := '0'; 
signal C_31_S_5_L_5_out : std_logic := '0'; 
signal C_32_S_0_L_0_out : std_logic := '0'; 
signal C_32_S_0_L_1_out : std_logic := '0'; 
signal C_32_S_0_L_2_out : std_logic := '0'; 
signal C_32_S_0_L_3_out : std_logic := '0'; 
signal C_32_S_0_L_4_out : std_logic := '0'; 
signal C_32_S_0_L_5_out : std_logic := '0'; 
signal C_32_S_1_L_0_out : std_logic := '0'; 
signal C_32_S_1_L_1_out : std_logic := '0'; 
signal C_32_S_1_L_2_out : std_logic := '0'; 
signal C_32_S_1_L_3_out : std_logic := '0'; 
signal C_32_S_1_L_4_out : std_logic := '0'; 
signal C_32_S_1_L_5_out : std_logic := '0'; 
signal C_32_S_2_L_0_out : std_logic := '0'; 
signal C_32_S_2_L_1_out : std_logic := '0'; 
signal C_32_S_2_L_2_out : std_logic := '0'; 
signal C_32_S_2_L_3_out : std_logic := '0'; 
signal C_32_S_2_L_4_out : std_logic := '0'; 
signal C_32_S_2_L_5_out : std_logic := '0'; 
signal C_32_S_3_L_0_out : std_logic := '0'; 
signal C_32_S_3_L_1_out : std_logic := '0'; 
signal C_32_S_3_L_2_out : std_logic := '0'; 
signal C_32_S_3_L_3_out : std_logic := '0'; 
signal C_32_S_3_L_4_out : std_logic := '0'; 
signal C_32_S_3_L_5_out : std_logic := '0'; 
signal C_32_S_4_L_0_out : std_logic := '0'; 
signal C_32_S_4_L_1_out : std_logic := '0'; 
signal C_32_S_4_L_2_out : std_logic := '0'; 
signal C_32_S_4_L_3_out : std_logic := '0'; 
signal C_32_S_4_L_4_out : std_logic := '0'; 
signal C_32_S_4_L_5_out : std_logic := '0'; 
signal C_32_S_5_L_0_out : std_logic := '0'; 
signal C_32_S_5_L_1_out : std_logic := '0'; 
signal C_32_S_5_L_2_out : std_logic := '0'; 
signal C_32_S_5_L_3_out : std_logic := '0'; 
signal C_32_S_5_L_4_out : std_logic := '0'; 
signal C_32_S_5_L_5_out : std_logic := '0'; 
signal C_33_S_0_L_0_out : std_logic := '0'; 
signal C_33_S_0_L_1_out : std_logic := '0'; 
signal C_33_S_0_L_2_out : std_logic := '0'; 
signal C_33_S_0_L_3_out : std_logic := '0'; 
signal C_33_S_0_L_4_out : std_logic := '0'; 
signal C_33_S_0_L_5_out : std_logic := '0'; 
signal C_33_S_1_L_0_out : std_logic := '0'; 
signal C_33_S_1_L_1_out : std_logic := '0'; 
signal C_33_S_1_L_2_out : std_logic := '0'; 
signal C_33_S_1_L_3_out : std_logic := '0'; 
signal C_33_S_1_L_4_out : std_logic := '0'; 
signal C_33_S_1_L_5_out : std_logic := '0'; 
signal C_33_S_2_L_0_out : std_logic := '0'; 
signal C_33_S_2_L_1_out : std_logic := '0'; 
signal C_33_S_2_L_2_out : std_logic := '0'; 
signal C_33_S_2_L_3_out : std_logic := '0'; 
signal C_33_S_2_L_4_out : std_logic := '0'; 
signal C_33_S_2_L_5_out : std_logic := '0'; 
signal C_33_S_3_L_0_out : std_logic := '0'; 
signal C_33_S_3_L_1_out : std_logic := '0'; 
signal C_33_S_3_L_2_out : std_logic := '0'; 
signal C_33_S_3_L_3_out : std_logic := '0'; 
signal C_33_S_3_L_4_out : std_logic := '0'; 
signal C_33_S_3_L_5_out : std_logic := '0'; 
signal C_33_S_4_L_0_out : std_logic := '0'; 
signal C_33_S_4_L_1_out : std_logic := '0'; 
signal C_33_S_4_L_2_out : std_logic := '0'; 
signal C_33_S_4_L_3_out : std_logic := '0'; 
signal C_33_S_4_L_4_out : std_logic := '0'; 
signal C_33_S_4_L_5_out : std_logic := '0'; 
signal C_33_S_5_L_0_out : std_logic := '0'; 
signal C_33_S_5_L_1_out : std_logic := '0'; 
signal C_33_S_5_L_2_out : std_logic := '0'; 
signal C_33_S_5_L_3_out : std_logic := '0'; 
signal C_33_S_5_L_4_out : std_logic := '0'; 
signal C_33_S_5_L_5_out : std_logic := '0'; 
signal C_34_S_0_L_0_out : std_logic := '0'; 
signal C_34_S_0_L_1_out : std_logic := '0'; 
signal C_34_S_0_L_2_out : std_logic := '0'; 
signal C_34_S_0_L_3_out : std_logic := '0'; 
signal C_34_S_0_L_4_out : std_logic := '0'; 
signal C_34_S_0_L_5_out : std_logic := '0'; 
signal C_34_S_1_L_0_out : std_logic := '0'; 
signal C_34_S_1_L_1_out : std_logic := '0'; 
signal C_34_S_1_L_2_out : std_logic := '0'; 
signal C_34_S_1_L_3_out : std_logic := '0'; 
signal C_34_S_1_L_4_out : std_logic := '0'; 
signal C_34_S_1_L_5_out : std_logic := '0'; 
signal C_34_S_2_L_0_out : std_logic := '0'; 
signal C_34_S_2_L_1_out : std_logic := '0'; 
signal C_34_S_2_L_2_out : std_logic := '0'; 
signal C_34_S_2_L_3_out : std_logic := '0'; 
signal C_34_S_2_L_4_out : std_logic := '0'; 
signal C_34_S_2_L_5_out : std_logic := '0'; 
signal C_34_S_3_L_0_out : std_logic := '0'; 
signal C_34_S_3_L_1_out : std_logic := '0'; 
signal C_34_S_3_L_2_out : std_logic := '0'; 
signal C_34_S_3_L_3_out : std_logic := '0'; 
signal C_34_S_3_L_4_out : std_logic := '0'; 
signal C_34_S_3_L_5_out : std_logic := '0'; 
signal C_34_S_4_L_0_out : std_logic := '0'; 
signal C_34_S_4_L_1_out : std_logic := '0'; 
signal C_34_S_4_L_2_out : std_logic := '0'; 
signal C_34_S_4_L_3_out : std_logic := '0'; 
signal C_34_S_4_L_4_out : std_logic := '0'; 
signal C_34_S_4_L_5_out : std_logic := '0'; 
signal C_34_S_5_L_0_out : std_logic := '0'; 
signal C_34_S_5_L_1_out : std_logic := '0'; 
signal C_34_S_5_L_2_out : std_logic := '0'; 
signal C_34_S_5_L_3_out : std_logic := '0'; 
signal C_34_S_5_L_4_out : std_logic := '0'; 
signal C_34_S_5_L_5_out : std_logic := '0'; 
signal C_35_S_0_L_0_out : std_logic := '0'; 
signal C_35_S_0_L_1_out : std_logic := '0'; 
signal C_35_S_0_L_2_out : std_logic := '0'; 
signal C_35_S_0_L_3_out : std_logic := '0'; 
signal C_35_S_0_L_4_out : std_logic := '0'; 
signal C_35_S_0_L_5_out : std_logic := '0'; 
signal C_35_S_1_L_0_out : std_logic := '0'; 
signal C_35_S_1_L_1_out : std_logic := '0'; 
signal C_35_S_1_L_2_out : std_logic := '0'; 
signal C_35_S_1_L_3_out : std_logic := '0'; 
signal C_35_S_1_L_4_out : std_logic := '0'; 
signal C_35_S_1_L_5_out : std_logic := '0'; 
signal C_35_S_2_L_0_out : std_logic := '0'; 
signal C_35_S_2_L_1_out : std_logic := '0'; 
signal C_35_S_2_L_2_out : std_logic := '0'; 
signal C_35_S_2_L_3_out : std_logic := '0'; 
signal C_35_S_2_L_4_out : std_logic := '0'; 
signal C_35_S_2_L_5_out : std_logic := '0'; 
signal C_35_S_3_L_0_out : std_logic := '0'; 
signal C_35_S_3_L_1_out : std_logic := '0'; 
signal C_35_S_3_L_2_out : std_logic := '0'; 
signal C_35_S_3_L_3_out : std_logic := '0'; 
signal C_35_S_3_L_4_out : std_logic := '0'; 
signal C_35_S_3_L_5_out : std_logic := '0'; 
signal C_35_S_4_L_0_out : std_logic := '0'; 
signal C_35_S_4_L_1_out : std_logic := '0'; 
signal C_35_S_4_L_2_out : std_logic := '0'; 
signal C_35_S_4_L_3_out : std_logic := '0'; 
signal C_35_S_4_L_4_out : std_logic := '0'; 
signal C_35_S_4_L_5_out : std_logic := '0'; 
signal C_35_S_5_L_0_out : std_logic := '0'; 
signal C_35_S_5_L_1_out : std_logic := '0'; 
signal C_35_S_5_L_2_out : std_logic := '0'; 
signal C_35_S_5_L_3_out : std_logic := '0'; 
signal C_35_S_5_L_4_out : std_logic := '0'; 
signal C_35_S_5_L_5_out : std_logic := '0'; 
signal C_36_S_0_L_0_out : std_logic := '0'; 
signal C_36_S_0_L_1_out : std_logic := '0'; 
signal C_36_S_0_L_2_out : std_logic := '0'; 
signal C_36_S_0_L_3_out : std_logic := '0'; 
signal C_36_S_0_L_4_out : std_logic := '0'; 
signal C_36_S_0_L_5_out : std_logic := '0'; 
signal C_36_S_1_L_0_out : std_logic := '0'; 
signal C_36_S_1_L_1_out : std_logic := '0'; 
signal C_36_S_1_L_2_out : std_logic := '0'; 
signal C_36_S_1_L_3_out : std_logic := '0'; 
signal C_36_S_1_L_4_out : std_logic := '0'; 
signal C_36_S_1_L_5_out : std_logic := '0'; 
signal C_36_S_2_L_0_out : std_logic := '0'; 
signal C_36_S_2_L_1_out : std_logic := '0'; 
signal C_36_S_2_L_2_out : std_logic := '0'; 
signal C_36_S_2_L_3_out : std_logic := '0'; 
signal C_36_S_2_L_4_out : std_logic := '0'; 
signal C_36_S_2_L_5_out : std_logic := '0'; 
signal C_36_S_3_L_0_out : std_logic := '0'; 
signal C_36_S_3_L_1_out : std_logic := '0'; 
signal C_36_S_3_L_2_out : std_logic := '0'; 
signal C_36_S_3_L_3_out : std_logic := '0'; 
signal C_36_S_3_L_4_out : std_logic := '0'; 
signal C_36_S_3_L_5_out : std_logic := '0'; 
signal C_36_S_4_L_0_out : std_logic := '0'; 
signal C_36_S_4_L_1_out : std_logic := '0'; 
signal C_36_S_4_L_2_out : std_logic := '0'; 
signal C_36_S_4_L_3_out : std_logic := '0'; 
signal C_36_S_4_L_4_out : std_logic := '0'; 
signal C_36_S_4_L_5_out : std_logic := '0'; 
signal C_36_S_5_L_0_out : std_logic := '0'; 
signal C_36_S_5_L_1_out : std_logic := '0'; 
signal C_36_S_5_L_2_out : std_logic := '0'; 
signal C_36_S_5_L_3_out : std_logic := '0'; 
signal C_36_S_5_L_4_out : std_logic := '0'; 
signal C_36_S_5_L_5_out : std_logic := '0'; 
signal C_37_S_0_L_0_out : std_logic := '0'; 
signal C_37_S_0_L_1_out : std_logic := '0'; 
signal C_37_S_0_L_2_out : std_logic := '0'; 
signal C_37_S_0_L_3_out : std_logic := '0'; 
signal C_37_S_0_L_4_out : std_logic := '0'; 
signal C_37_S_0_L_5_out : std_logic := '0'; 
signal C_37_S_1_L_0_out : std_logic := '0'; 
signal C_37_S_1_L_1_out : std_logic := '0'; 
signal C_37_S_1_L_2_out : std_logic := '0'; 
signal C_37_S_1_L_3_out : std_logic := '0'; 
signal C_37_S_1_L_4_out : std_logic := '0'; 
signal C_37_S_1_L_5_out : std_logic := '0'; 
signal C_37_S_2_L_0_out : std_logic := '0'; 
signal C_37_S_2_L_1_out : std_logic := '0'; 
signal C_37_S_2_L_2_out : std_logic := '0'; 
signal C_37_S_2_L_3_out : std_logic := '0'; 
signal C_37_S_2_L_4_out : std_logic := '0'; 
signal C_37_S_2_L_5_out : std_logic := '0'; 
signal C_37_S_3_L_0_out : std_logic := '0'; 
signal C_37_S_3_L_1_out : std_logic := '0'; 
signal C_37_S_3_L_2_out : std_logic := '0'; 
signal C_37_S_3_L_3_out : std_logic := '0'; 
signal C_37_S_3_L_4_out : std_logic := '0'; 
signal C_37_S_3_L_5_out : std_logic := '0'; 
signal C_37_S_4_L_0_out : std_logic := '0'; 
signal C_37_S_4_L_1_out : std_logic := '0'; 
signal C_37_S_4_L_2_out : std_logic := '0'; 
signal C_37_S_4_L_3_out : std_logic := '0'; 
signal C_37_S_4_L_4_out : std_logic := '0'; 
signal C_37_S_4_L_5_out : std_logic := '0'; 
signal C_37_S_5_L_0_out : std_logic := '0'; 
signal C_37_S_5_L_1_out : std_logic := '0'; 
signal C_37_S_5_L_2_out : std_logic := '0'; 
signal C_37_S_5_L_3_out : std_logic := '0'; 
signal C_37_S_5_L_4_out : std_logic := '0'; 
signal C_37_S_5_L_5_out : std_logic := '0'; 
signal C_38_S_0_L_0_out : std_logic := '0'; 
signal C_38_S_0_L_1_out : std_logic := '0'; 
signal C_38_S_0_L_2_out : std_logic := '0'; 
signal C_38_S_0_L_3_out : std_logic := '0'; 
signal C_38_S_0_L_4_out : std_logic := '0'; 
signal C_38_S_0_L_5_out : std_logic := '0'; 
signal C_38_S_1_L_0_out : std_logic := '0'; 
signal C_38_S_1_L_1_out : std_logic := '0'; 
signal C_38_S_1_L_2_out : std_logic := '0'; 
signal C_38_S_1_L_3_out : std_logic := '0'; 
signal C_38_S_1_L_4_out : std_logic := '0'; 
signal C_38_S_1_L_5_out : std_logic := '0'; 
signal C_38_S_2_L_0_out : std_logic := '0'; 
signal C_38_S_2_L_1_out : std_logic := '0'; 
signal C_38_S_2_L_2_out : std_logic := '0'; 
signal C_38_S_2_L_3_out : std_logic := '0'; 
signal C_38_S_2_L_4_out : std_logic := '0'; 
signal C_38_S_2_L_5_out : std_logic := '0'; 
signal C_38_S_3_L_0_out : std_logic := '0'; 
signal C_38_S_3_L_1_out : std_logic := '0'; 
signal C_38_S_3_L_2_out : std_logic := '0'; 
signal C_38_S_3_L_3_out : std_logic := '0'; 
signal C_38_S_3_L_4_out : std_logic := '0'; 
signal C_38_S_3_L_5_out : std_logic := '0'; 
signal C_38_S_4_L_0_out : std_logic := '0'; 
signal C_38_S_4_L_1_out : std_logic := '0'; 
signal C_38_S_4_L_2_out : std_logic := '0'; 
signal C_38_S_4_L_3_out : std_logic := '0'; 
signal C_38_S_4_L_4_out : std_logic := '0'; 
signal C_38_S_4_L_5_out : std_logic := '0'; 
signal C_38_S_5_L_0_out : std_logic := '0'; 
signal C_38_S_5_L_1_out : std_logic := '0'; 
signal C_38_S_5_L_2_out : std_logic := '0'; 
signal C_38_S_5_L_3_out : std_logic := '0'; 
signal C_38_S_5_L_4_out : std_logic := '0'; 
signal C_38_S_5_L_5_out : std_logic := '0'; 
signal C_39_S_0_L_0_out : std_logic := '0'; 
signal C_39_S_0_L_1_out : std_logic := '0'; 
signal C_39_S_0_L_2_out : std_logic := '0'; 
signal C_39_S_0_L_3_out : std_logic := '0'; 
signal C_39_S_0_L_4_out : std_logic := '0'; 
signal C_39_S_0_L_5_out : std_logic := '0'; 
signal C_39_S_1_L_0_out : std_logic := '0'; 
signal C_39_S_1_L_1_out : std_logic := '0'; 
signal C_39_S_1_L_2_out : std_logic := '0'; 
signal C_39_S_1_L_3_out : std_logic := '0'; 
signal C_39_S_1_L_4_out : std_logic := '0'; 
signal C_39_S_1_L_5_out : std_logic := '0'; 
signal C_39_S_2_L_0_out : std_logic := '0'; 
signal C_39_S_2_L_1_out : std_logic := '0'; 
signal C_39_S_2_L_2_out : std_logic := '0'; 
signal C_39_S_2_L_3_out : std_logic := '0'; 
signal C_39_S_2_L_4_out : std_logic := '0'; 
signal C_39_S_2_L_5_out : std_logic := '0'; 
signal C_39_S_3_L_0_out : std_logic := '0'; 
signal C_39_S_3_L_1_out : std_logic := '0'; 
signal C_39_S_3_L_2_out : std_logic := '0'; 
signal C_39_S_3_L_3_out : std_logic := '0'; 
signal C_39_S_3_L_4_out : std_logic := '0'; 
signal C_39_S_3_L_5_out : std_logic := '0'; 
signal C_39_S_4_L_0_out : std_logic := '0'; 
signal C_39_S_4_L_1_out : std_logic := '0'; 
signal C_39_S_4_L_2_out : std_logic := '0'; 
signal C_39_S_4_L_3_out : std_logic := '0'; 
signal C_39_S_4_L_4_out : std_logic := '0'; 
signal C_39_S_4_L_5_out : std_logic := '0'; 
signal C_39_S_5_L_0_out : std_logic := '0'; 
signal C_39_S_5_L_1_out : std_logic := '0'; 
signal C_39_S_5_L_2_out : std_logic := '0'; 
signal C_39_S_5_L_3_out : std_logic := '0'; 
signal C_39_S_5_L_4_out : std_logic := '0'; 
signal C_39_S_5_L_5_out : std_logic := '0'; 
signal C_40_S_0_L_0_out : std_logic := '0'; 
signal C_40_S_0_L_1_out : std_logic := '0'; 
signal C_40_S_0_L_2_out : std_logic := '0'; 
signal C_40_S_0_L_3_out : std_logic := '0'; 
signal C_40_S_0_L_4_out : std_logic := '0'; 
signal C_40_S_0_L_5_out : std_logic := '0'; 
signal C_40_S_1_L_0_out : std_logic := '0'; 
signal C_40_S_1_L_1_out : std_logic := '0'; 
signal C_40_S_1_L_2_out : std_logic := '0'; 
signal C_40_S_1_L_3_out : std_logic := '0'; 
signal C_40_S_1_L_4_out : std_logic := '0'; 
signal C_40_S_1_L_5_out : std_logic := '0'; 
signal C_40_S_2_L_0_out : std_logic := '0'; 
signal C_40_S_2_L_1_out : std_logic := '0'; 
signal C_40_S_2_L_2_out : std_logic := '0'; 
signal C_40_S_2_L_3_out : std_logic := '0'; 
signal C_40_S_2_L_4_out : std_logic := '0'; 
signal C_40_S_2_L_5_out : std_logic := '0'; 
signal C_40_S_3_L_0_out : std_logic := '0'; 
signal C_40_S_3_L_1_out : std_logic := '0'; 
signal C_40_S_3_L_2_out : std_logic := '0'; 
signal C_40_S_3_L_3_out : std_logic := '0'; 
signal C_40_S_3_L_4_out : std_logic := '0'; 
signal C_40_S_3_L_5_out : std_logic := '0'; 
signal C_40_S_4_L_0_out : std_logic := '0'; 
signal C_40_S_4_L_1_out : std_logic := '0'; 
signal C_40_S_4_L_2_out : std_logic := '0'; 
signal C_40_S_4_L_3_out : std_logic := '0'; 
signal C_40_S_4_L_4_out : std_logic := '0'; 
signal C_40_S_4_L_5_out : std_logic := '0'; 
signal C_40_S_5_L_0_out : std_logic := '0'; 
signal C_40_S_5_L_1_out : std_logic := '0'; 
signal C_40_S_5_L_2_out : std_logic := '0'; 
signal C_40_S_5_L_3_out : std_logic := '0'; 
signal C_40_S_5_L_4_out : std_logic := '0'; 
signal C_40_S_5_L_5_out : std_logic := '0'; 
signal C_41_S_0_L_0_out : std_logic := '0'; 
signal C_41_S_0_L_1_out : std_logic := '0'; 
signal C_41_S_0_L_2_out : std_logic := '0'; 
signal C_41_S_0_L_3_out : std_logic := '0'; 
signal C_41_S_0_L_4_out : std_logic := '0'; 
signal C_41_S_0_L_5_out : std_logic := '0'; 
signal C_41_S_1_L_0_out : std_logic := '0'; 
signal C_41_S_1_L_1_out : std_logic := '0'; 
signal C_41_S_1_L_2_out : std_logic := '0'; 
signal C_41_S_1_L_3_out : std_logic := '0'; 
signal C_41_S_1_L_4_out : std_logic := '0'; 
signal C_41_S_1_L_5_out : std_logic := '0'; 
signal C_41_S_2_L_0_out : std_logic := '0'; 
signal C_41_S_2_L_1_out : std_logic := '0'; 
signal C_41_S_2_L_2_out : std_logic := '0'; 
signal C_41_S_2_L_3_out : std_logic := '0'; 
signal C_41_S_2_L_4_out : std_logic := '0'; 
signal C_41_S_2_L_5_out : std_logic := '0'; 
signal C_41_S_3_L_0_out : std_logic := '0'; 
signal C_41_S_3_L_1_out : std_logic := '0'; 
signal C_41_S_3_L_2_out : std_logic := '0'; 
signal C_41_S_3_L_3_out : std_logic := '0'; 
signal C_41_S_3_L_4_out : std_logic := '0'; 
signal C_41_S_3_L_5_out : std_logic := '0'; 
signal C_41_S_4_L_0_out : std_logic := '0'; 
signal C_41_S_4_L_1_out : std_logic := '0'; 
signal C_41_S_4_L_2_out : std_logic := '0'; 
signal C_41_S_4_L_3_out : std_logic := '0'; 
signal C_41_S_4_L_4_out : std_logic := '0'; 
signal C_41_S_4_L_5_out : std_logic := '0'; 
signal C_41_S_5_L_0_out : std_logic := '0'; 
signal C_41_S_5_L_1_out : std_logic := '0'; 
signal C_41_S_5_L_2_out : std_logic := '0'; 
signal C_41_S_5_L_3_out : std_logic := '0'; 
signal C_41_S_5_L_4_out : std_logic := '0'; 
signal C_41_S_5_L_5_out : std_logic := '0'; 
signal C_42_S_0_L_0_out : std_logic := '0'; 
signal C_42_S_0_L_1_out : std_logic := '0'; 
signal C_42_S_0_L_2_out : std_logic := '0'; 
signal C_42_S_0_L_3_out : std_logic := '0'; 
signal C_42_S_0_L_4_out : std_logic := '0'; 
signal C_42_S_0_L_5_out : std_logic := '0'; 
signal C_42_S_1_L_0_out : std_logic := '0'; 
signal C_42_S_1_L_1_out : std_logic := '0'; 
signal C_42_S_1_L_2_out : std_logic := '0'; 
signal C_42_S_1_L_3_out : std_logic := '0'; 
signal C_42_S_1_L_4_out : std_logic := '0'; 
signal C_42_S_1_L_5_out : std_logic := '0'; 
signal C_42_S_2_L_0_out : std_logic := '0'; 
signal C_42_S_2_L_1_out : std_logic := '0'; 
signal C_42_S_2_L_2_out : std_logic := '0'; 
signal C_42_S_2_L_3_out : std_logic := '0'; 
signal C_42_S_2_L_4_out : std_logic := '0'; 
signal C_42_S_2_L_5_out : std_logic := '0'; 
signal C_42_S_3_L_0_out : std_logic := '0'; 
signal C_42_S_3_L_1_out : std_logic := '0'; 
signal C_42_S_3_L_2_out : std_logic := '0'; 
signal C_42_S_3_L_3_out : std_logic := '0'; 
signal C_42_S_3_L_4_out : std_logic := '0'; 
signal C_42_S_3_L_5_out : std_logic := '0'; 
signal C_42_S_4_L_0_out : std_logic := '0'; 
signal C_42_S_4_L_1_out : std_logic := '0'; 
signal C_42_S_4_L_2_out : std_logic := '0'; 
signal C_42_S_4_L_3_out : std_logic := '0'; 
signal C_42_S_4_L_4_out : std_logic := '0'; 
signal C_42_S_4_L_5_out : std_logic := '0'; 
signal C_42_S_5_L_0_out : std_logic := '0'; 
signal C_42_S_5_L_1_out : std_logic := '0'; 
signal C_42_S_5_L_2_out : std_logic := '0'; 
signal C_42_S_5_L_3_out : std_logic := '0'; 
signal C_42_S_5_L_4_out : std_logic := '0'; 
signal C_42_S_5_L_5_out : std_logic := '0'; 
signal C_43_S_0_L_0_out : std_logic := '0'; 
signal C_43_S_0_L_1_out : std_logic := '0'; 
signal C_43_S_0_L_2_out : std_logic := '0'; 
signal C_43_S_0_L_3_out : std_logic := '0'; 
signal C_43_S_0_L_4_out : std_logic := '0'; 
signal C_43_S_0_L_5_out : std_logic := '0'; 
signal C_43_S_1_L_0_out : std_logic := '0'; 
signal C_43_S_1_L_1_out : std_logic := '0'; 
signal C_43_S_1_L_2_out : std_logic := '0'; 
signal C_43_S_1_L_3_out : std_logic := '0'; 
signal C_43_S_1_L_4_out : std_logic := '0'; 
signal C_43_S_1_L_5_out : std_logic := '0'; 
signal C_43_S_2_L_0_out : std_logic := '0'; 
signal C_43_S_2_L_1_out : std_logic := '0'; 
signal C_43_S_2_L_2_out : std_logic := '0'; 
signal C_43_S_2_L_3_out : std_logic := '0'; 
signal C_43_S_2_L_4_out : std_logic := '0'; 
signal C_43_S_2_L_5_out : std_logic := '0'; 
signal C_43_S_3_L_0_out : std_logic := '0'; 
signal C_43_S_3_L_1_out : std_logic := '0'; 
signal C_43_S_3_L_2_out : std_logic := '0'; 
signal C_43_S_3_L_3_out : std_logic := '0'; 
signal C_43_S_3_L_4_out : std_logic := '0'; 
signal C_43_S_3_L_5_out : std_logic := '0'; 
signal C_43_S_4_L_0_out : std_logic := '0'; 
signal C_43_S_4_L_1_out : std_logic := '0'; 
signal C_43_S_4_L_2_out : std_logic := '0'; 
signal C_43_S_4_L_3_out : std_logic := '0'; 
signal C_43_S_4_L_4_out : std_logic := '0'; 
signal C_43_S_4_L_5_out : std_logic := '0'; 
signal C_43_S_5_L_0_out : std_logic := '0'; 
signal C_43_S_5_L_1_out : std_logic := '0'; 
signal C_43_S_5_L_2_out : std_logic := '0'; 
signal C_43_S_5_L_3_out : std_logic := '0'; 
signal C_43_S_5_L_4_out : std_logic := '0'; 
signal C_43_S_5_L_5_out : std_logic := '0'; 
signal C_44_S_0_L_0_out : std_logic := '0'; 
signal C_44_S_0_L_1_out : std_logic := '0'; 
signal C_44_S_0_L_2_out : std_logic := '0'; 
signal C_44_S_0_L_3_out : std_logic := '0'; 
signal C_44_S_0_L_4_out : std_logic := '0'; 
signal C_44_S_0_L_5_out : std_logic := '0'; 
signal C_44_S_1_L_0_out : std_logic := '0'; 
signal C_44_S_1_L_1_out : std_logic := '0'; 
signal C_44_S_1_L_2_out : std_logic := '0'; 
signal C_44_S_1_L_3_out : std_logic := '0'; 
signal C_44_S_1_L_4_out : std_logic := '0'; 
signal C_44_S_1_L_5_out : std_logic := '0'; 
signal C_44_S_2_L_0_out : std_logic := '0'; 
signal C_44_S_2_L_1_out : std_logic := '0'; 
signal C_44_S_2_L_2_out : std_logic := '0'; 
signal C_44_S_2_L_3_out : std_logic := '0'; 
signal C_44_S_2_L_4_out : std_logic := '0'; 
signal C_44_S_2_L_5_out : std_logic := '0'; 
signal C_44_S_3_L_0_out : std_logic := '0'; 
signal C_44_S_3_L_1_out : std_logic := '0'; 
signal C_44_S_3_L_2_out : std_logic := '0'; 
signal C_44_S_3_L_3_out : std_logic := '0'; 
signal C_44_S_3_L_4_out : std_logic := '0'; 
signal C_44_S_3_L_5_out : std_logic := '0'; 
signal C_44_S_4_L_0_out : std_logic := '0'; 
signal C_44_S_4_L_1_out : std_logic := '0'; 
signal C_44_S_4_L_2_out : std_logic := '0'; 
signal C_44_S_4_L_3_out : std_logic := '0'; 
signal C_44_S_4_L_4_out : std_logic := '0'; 
signal C_44_S_4_L_5_out : std_logic := '0'; 
signal C_44_S_5_L_0_out : std_logic := '0'; 
signal C_44_S_5_L_1_out : std_logic := '0'; 
signal C_44_S_5_L_2_out : std_logic := '0'; 
signal C_44_S_5_L_3_out : std_logic := '0'; 
signal C_44_S_5_L_4_out : std_logic := '0'; 
signal C_44_S_5_L_5_out : std_logic := '0'; 
signal C_45_S_0_L_0_out : std_logic := '0'; 
signal C_45_S_0_L_1_out : std_logic := '0'; 
signal C_45_S_0_L_2_out : std_logic := '0'; 
signal C_45_S_0_L_3_out : std_logic := '0'; 
signal C_45_S_0_L_4_out : std_logic := '0'; 
signal C_45_S_0_L_5_out : std_logic := '0'; 
signal C_45_S_1_L_0_out : std_logic := '0'; 
signal C_45_S_1_L_1_out : std_logic := '0'; 
signal C_45_S_1_L_2_out : std_logic := '0'; 
signal C_45_S_1_L_3_out : std_logic := '0'; 
signal C_45_S_1_L_4_out : std_logic := '0'; 
signal C_45_S_1_L_5_out : std_logic := '0'; 
signal C_45_S_2_L_0_out : std_logic := '0'; 
signal C_45_S_2_L_1_out : std_logic := '0'; 
signal C_45_S_2_L_2_out : std_logic := '0'; 
signal C_45_S_2_L_3_out : std_logic := '0'; 
signal C_45_S_2_L_4_out : std_logic := '0'; 
signal C_45_S_2_L_5_out : std_logic := '0'; 
signal C_45_S_3_L_0_out : std_logic := '0'; 
signal C_45_S_3_L_1_out : std_logic := '0'; 
signal C_45_S_3_L_2_out : std_logic := '0'; 
signal C_45_S_3_L_3_out : std_logic := '0'; 
signal C_45_S_3_L_4_out : std_logic := '0'; 
signal C_45_S_3_L_5_out : std_logic := '0'; 
signal C_45_S_4_L_0_out : std_logic := '0'; 
signal C_45_S_4_L_1_out : std_logic := '0'; 
signal C_45_S_4_L_2_out : std_logic := '0'; 
signal C_45_S_4_L_3_out : std_logic := '0'; 
signal C_45_S_4_L_4_out : std_logic := '0'; 
signal C_45_S_4_L_5_out : std_logic := '0'; 
signal C_45_S_5_L_0_out : std_logic := '0'; 
signal C_45_S_5_L_1_out : std_logic := '0'; 
signal C_45_S_5_L_2_out : std_logic := '0'; 
signal C_45_S_5_L_3_out : std_logic := '0'; 
signal C_45_S_5_L_4_out : std_logic := '0'; 
signal C_45_S_5_L_5_out : std_logic := '0'; 
signal C_46_S_0_L_0_out : std_logic := '0'; 
signal C_46_S_0_L_1_out : std_logic := '0'; 
signal C_46_S_0_L_2_out : std_logic := '0'; 
signal C_46_S_0_L_3_out : std_logic := '0'; 
signal C_46_S_0_L_4_out : std_logic := '0'; 
signal C_46_S_0_L_5_out : std_logic := '0'; 
signal C_46_S_1_L_0_out : std_logic := '0'; 
signal C_46_S_1_L_1_out : std_logic := '0'; 
signal C_46_S_1_L_2_out : std_logic := '0'; 
signal C_46_S_1_L_3_out : std_logic := '0'; 
signal C_46_S_1_L_4_out : std_logic := '0'; 
signal C_46_S_1_L_5_out : std_logic := '0'; 
signal C_46_S_2_L_0_out : std_logic := '0'; 
signal C_46_S_2_L_1_out : std_logic := '0'; 
signal C_46_S_2_L_2_out : std_logic := '0'; 
signal C_46_S_2_L_3_out : std_logic := '0'; 
signal C_46_S_2_L_4_out : std_logic := '0'; 
signal C_46_S_2_L_5_out : std_logic := '0'; 
signal C_46_S_3_L_0_out : std_logic := '0'; 
signal C_46_S_3_L_1_out : std_logic := '0'; 
signal C_46_S_3_L_2_out : std_logic := '0'; 
signal C_46_S_3_L_3_out : std_logic := '0'; 
signal C_46_S_3_L_4_out : std_logic := '0'; 
signal C_46_S_3_L_5_out : std_logic := '0'; 
signal C_46_S_4_L_0_out : std_logic := '0'; 
signal C_46_S_4_L_1_out : std_logic := '0'; 
signal C_46_S_4_L_2_out : std_logic := '0'; 
signal C_46_S_4_L_3_out : std_logic := '0'; 
signal C_46_S_4_L_4_out : std_logic := '0'; 
signal C_46_S_4_L_5_out : std_logic := '0'; 
signal C_46_S_5_L_0_out : std_logic := '0'; 
signal C_46_S_5_L_1_out : std_logic := '0'; 
signal C_46_S_5_L_2_out : std_logic := '0'; 
signal C_46_S_5_L_3_out : std_logic := '0'; 
signal C_46_S_5_L_4_out : std_logic := '0'; 
signal C_46_S_5_L_5_out : std_logic := '0'; 
signal C_47_S_0_L_0_out : std_logic := '0'; 
signal C_47_S_0_L_1_out : std_logic := '0'; 
signal C_47_S_0_L_2_out : std_logic := '0'; 
signal C_47_S_0_L_3_out : std_logic := '0'; 
signal C_47_S_0_L_4_out : std_logic := '0'; 
signal C_47_S_0_L_5_out : std_logic := '0'; 
signal C_47_S_1_L_0_out : std_logic := '0'; 
signal C_47_S_1_L_1_out : std_logic := '0'; 
signal C_47_S_1_L_2_out : std_logic := '0'; 
signal C_47_S_1_L_3_out : std_logic := '0'; 
signal C_47_S_1_L_4_out : std_logic := '0'; 
signal C_47_S_1_L_5_out : std_logic := '0'; 
signal C_47_S_2_L_0_out : std_logic := '0'; 
signal C_47_S_2_L_1_out : std_logic := '0'; 
signal C_47_S_2_L_2_out : std_logic := '0'; 
signal C_47_S_2_L_3_out : std_logic := '0'; 
signal C_47_S_2_L_4_out : std_logic := '0'; 
signal C_47_S_2_L_5_out : std_logic := '0'; 
signal C_47_S_3_L_0_out : std_logic := '0'; 
signal C_47_S_3_L_1_out : std_logic := '0'; 
signal C_47_S_3_L_2_out : std_logic := '0'; 
signal C_47_S_3_L_3_out : std_logic := '0'; 
signal C_47_S_3_L_4_out : std_logic := '0'; 
signal C_47_S_3_L_5_out : std_logic := '0'; 
signal C_47_S_4_L_0_out : std_logic := '0'; 
signal C_47_S_4_L_1_out : std_logic := '0'; 
signal C_47_S_4_L_2_out : std_logic := '0'; 
signal C_47_S_4_L_3_out : std_logic := '0'; 
signal C_47_S_4_L_4_out : std_logic := '0'; 
signal C_47_S_4_L_5_out : std_logic := '0'; 
signal C_47_S_5_L_0_out : std_logic := '0'; 
signal C_47_S_5_L_1_out : std_logic := '0'; 
signal C_47_S_5_L_2_out : std_logic := '0'; 
signal C_47_S_5_L_3_out : std_logic := '0'; 
signal C_47_S_5_L_4_out : std_logic := '0'; 
signal C_47_S_5_L_5_out : std_logic := '0'; 
signal C_48_S_0_L_0_out : std_logic := '0'; 
signal C_48_S_0_L_1_out : std_logic := '0'; 
signal C_48_S_0_L_2_out : std_logic := '0'; 
signal C_48_S_0_L_3_out : std_logic := '0'; 
signal C_48_S_0_L_4_out : std_logic := '0'; 
signal C_48_S_0_L_5_out : std_logic := '0'; 
signal C_48_S_1_L_0_out : std_logic := '0'; 
signal C_48_S_1_L_1_out : std_logic := '0'; 
signal C_48_S_1_L_2_out : std_logic := '0'; 
signal C_48_S_1_L_3_out : std_logic := '0'; 
signal C_48_S_1_L_4_out : std_logic := '0'; 
signal C_48_S_1_L_5_out : std_logic := '0'; 
signal C_48_S_2_L_0_out : std_logic := '0'; 
signal C_48_S_2_L_1_out : std_logic := '0'; 
signal C_48_S_2_L_2_out : std_logic := '0'; 
signal C_48_S_2_L_3_out : std_logic := '0'; 
signal C_48_S_2_L_4_out : std_logic := '0'; 
signal C_48_S_2_L_5_out : std_logic := '0'; 
signal C_48_S_3_L_0_out : std_logic := '0'; 
signal C_48_S_3_L_1_out : std_logic := '0'; 
signal C_48_S_3_L_2_out : std_logic := '0'; 
signal C_48_S_3_L_3_out : std_logic := '0'; 
signal C_48_S_3_L_4_out : std_logic := '0'; 
signal C_48_S_3_L_5_out : std_logic := '0'; 
signal C_48_S_4_L_0_out : std_logic := '0'; 
signal C_48_S_4_L_1_out : std_logic := '0'; 
signal C_48_S_4_L_2_out : std_logic := '0'; 
signal C_48_S_4_L_3_out : std_logic := '0'; 
signal C_48_S_4_L_4_out : std_logic := '0'; 
signal C_48_S_4_L_5_out : std_logic := '0'; 
signal C_48_S_5_L_0_out : std_logic := '0'; 
signal C_48_S_5_L_1_out : std_logic := '0'; 
signal C_48_S_5_L_2_out : std_logic := '0'; 
signal C_48_S_5_L_3_out : std_logic := '0'; 
signal C_48_S_5_L_4_out : std_logic := '0'; 
signal C_48_S_5_L_5_out : std_logic := '0'; 
signal C_49_S_0_L_0_out : std_logic := '0'; 
signal C_49_S_0_L_1_out : std_logic := '0'; 
signal C_49_S_0_L_2_out : std_logic := '0'; 
signal C_49_S_0_L_3_out : std_logic := '0'; 
signal C_49_S_0_L_4_out : std_logic := '0'; 
signal C_49_S_0_L_5_out : std_logic := '0'; 
signal C_49_S_1_L_0_out : std_logic := '0'; 
signal C_49_S_1_L_1_out : std_logic := '0'; 
signal C_49_S_1_L_2_out : std_logic := '0'; 
signal C_49_S_1_L_3_out : std_logic := '0'; 
signal C_49_S_1_L_4_out : std_logic := '0'; 
signal C_49_S_1_L_5_out : std_logic := '0'; 
signal C_49_S_2_L_0_out : std_logic := '0'; 
signal C_49_S_2_L_1_out : std_logic := '0'; 
signal C_49_S_2_L_2_out : std_logic := '0'; 
signal C_49_S_2_L_3_out : std_logic := '0'; 
signal C_49_S_2_L_4_out : std_logic := '0'; 
signal C_49_S_2_L_5_out : std_logic := '0'; 
signal C_49_S_3_L_0_out : std_logic := '0'; 
signal C_49_S_3_L_1_out : std_logic := '0'; 
signal C_49_S_3_L_2_out : std_logic := '0'; 
signal C_49_S_3_L_3_out : std_logic := '0'; 
signal C_49_S_3_L_4_out : std_logic := '0'; 
signal C_49_S_3_L_5_out : std_logic := '0'; 
signal C_49_S_4_L_0_out : std_logic := '0'; 
signal C_49_S_4_L_1_out : std_logic := '0'; 
signal C_49_S_4_L_2_out : std_logic := '0'; 
signal C_49_S_4_L_3_out : std_logic := '0'; 
signal C_49_S_4_L_4_out : std_logic := '0'; 
signal C_49_S_4_L_5_out : std_logic := '0'; 
signal C_49_S_5_L_0_out : std_logic := '0'; 
signal C_49_S_5_L_1_out : std_logic := '0'; 
signal C_49_S_5_L_2_out : std_logic := '0'; 
signal C_49_S_5_L_3_out : std_logic := '0'; 
signal C_49_S_5_L_4_out : std_logic := '0'; 
signal C_49_S_5_L_5_out : std_logic := '0'; 
signal C_50_S_0_L_0_out : std_logic := '0'; 
signal C_50_S_0_L_1_out : std_logic := '0'; 
signal C_50_S_0_L_2_out : std_logic := '0'; 
signal C_50_S_0_L_3_out : std_logic := '0'; 
signal C_50_S_0_L_4_out : std_logic := '0'; 
signal C_50_S_0_L_5_out : std_logic := '0'; 
signal C_50_S_1_L_0_out : std_logic := '0'; 
signal C_50_S_1_L_1_out : std_logic := '0'; 
signal C_50_S_1_L_2_out : std_logic := '0'; 
signal C_50_S_1_L_3_out : std_logic := '0'; 
signal C_50_S_1_L_4_out : std_logic := '0'; 
signal C_50_S_1_L_5_out : std_logic := '0'; 
signal C_50_S_2_L_0_out : std_logic := '0'; 
signal C_50_S_2_L_1_out : std_logic := '0'; 
signal C_50_S_2_L_2_out : std_logic := '0'; 
signal C_50_S_2_L_3_out : std_logic := '0'; 
signal C_50_S_2_L_4_out : std_logic := '0'; 
signal C_50_S_2_L_5_out : std_logic := '0'; 
signal C_50_S_3_L_0_out : std_logic := '0'; 
signal C_50_S_3_L_1_out : std_logic := '0'; 
signal C_50_S_3_L_2_out : std_logic := '0'; 
signal C_50_S_3_L_3_out : std_logic := '0'; 
signal C_50_S_3_L_4_out : std_logic := '0'; 
signal C_50_S_3_L_5_out : std_logic := '0'; 
signal C_50_S_4_L_0_out : std_logic := '0'; 
signal C_50_S_4_L_1_out : std_logic := '0'; 
signal C_50_S_4_L_2_out : std_logic := '0'; 
signal C_50_S_4_L_3_out : std_logic := '0'; 
signal C_50_S_4_L_4_out : std_logic := '0'; 
signal C_50_S_4_L_5_out : std_logic := '0'; 
signal C_50_S_5_L_0_out : std_logic := '0'; 
signal C_50_S_5_L_1_out : std_logic := '0'; 
signal C_50_S_5_L_2_out : std_logic := '0'; 
signal C_50_S_5_L_3_out : std_logic := '0'; 
signal C_50_S_5_L_4_out : std_logic := '0'; 
signal C_50_S_5_L_5_out : std_logic := '0'; 
signal C_51_S_0_L_0_out : std_logic := '0'; 
signal C_51_S_0_L_1_out : std_logic := '0'; 
signal C_51_S_0_L_2_out : std_logic := '0'; 
signal C_51_S_0_L_3_out : std_logic := '0'; 
signal C_51_S_0_L_4_out : std_logic := '0'; 
signal C_51_S_0_L_5_out : std_logic := '0'; 
signal C_51_S_1_L_0_out : std_logic := '0'; 
signal C_51_S_1_L_1_out : std_logic := '0'; 
signal C_51_S_1_L_2_out : std_logic := '0'; 
signal C_51_S_1_L_3_out : std_logic := '0'; 
signal C_51_S_1_L_4_out : std_logic := '0'; 
signal C_51_S_1_L_5_out : std_logic := '0'; 
signal C_51_S_2_L_0_out : std_logic := '0'; 
signal C_51_S_2_L_1_out : std_logic := '0'; 
signal C_51_S_2_L_2_out : std_logic := '0'; 
signal C_51_S_2_L_3_out : std_logic := '0'; 
signal C_51_S_2_L_4_out : std_logic := '0'; 
signal C_51_S_2_L_5_out : std_logic := '0'; 
signal C_51_S_3_L_0_out : std_logic := '0'; 
signal C_51_S_3_L_1_out : std_logic := '0'; 
signal C_51_S_3_L_2_out : std_logic := '0'; 
signal C_51_S_3_L_3_out : std_logic := '0'; 
signal C_51_S_3_L_4_out : std_logic := '0'; 
signal C_51_S_3_L_5_out : std_logic := '0'; 
signal C_51_S_4_L_0_out : std_logic := '0'; 
signal C_51_S_4_L_1_out : std_logic := '0'; 
signal C_51_S_4_L_2_out : std_logic := '0'; 
signal C_51_S_4_L_3_out : std_logic := '0'; 
signal C_51_S_4_L_4_out : std_logic := '0'; 
signal C_51_S_4_L_5_out : std_logic := '0'; 
signal C_51_S_5_L_0_out : std_logic := '0'; 
signal C_51_S_5_L_1_out : std_logic := '0'; 
signal C_51_S_5_L_2_out : std_logic := '0'; 
signal C_51_S_5_L_3_out : std_logic := '0'; 
signal C_51_S_5_L_4_out : std_logic := '0'; 
signal C_51_S_5_L_5_out : std_logic := '0'; 
signal C_52_S_0_L_0_out : std_logic := '0'; 
signal C_52_S_0_L_1_out : std_logic := '0'; 
signal C_52_S_0_L_2_out : std_logic := '0'; 
signal C_52_S_0_L_3_out : std_logic := '0'; 
signal C_52_S_0_L_4_out : std_logic := '0'; 
signal C_52_S_0_L_5_out : std_logic := '0'; 
signal C_52_S_1_L_0_out : std_logic := '0'; 
signal C_52_S_1_L_1_out : std_logic := '0'; 
signal C_52_S_1_L_2_out : std_logic := '0'; 
signal C_52_S_1_L_3_out : std_logic := '0'; 
signal C_52_S_1_L_4_out : std_logic := '0'; 
signal C_52_S_1_L_5_out : std_logic := '0'; 
signal C_52_S_2_L_0_out : std_logic := '0'; 
signal C_52_S_2_L_1_out : std_logic := '0'; 
signal C_52_S_2_L_2_out : std_logic := '0'; 
signal C_52_S_2_L_3_out : std_logic := '0'; 
signal C_52_S_2_L_4_out : std_logic := '0'; 
signal C_52_S_2_L_5_out : std_logic := '0'; 
signal C_52_S_3_L_0_out : std_logic := '0'; 
signal C_52_S_3_L_1_out : std_logic := '0'; 
signal C_52_S_3_L_2_out : std_logic := '0'; 
signal C_52_S_3_L_3_out : std_logic := '0'; 
signal C_52_S_3_L_4_out : std_logic := '0'; 
signal C_52_S_3_L_5_out : std_logic := '0'; 
signal C_52_S_4_L_0_out : std_logic := '0'; 
signal C_52_S_4_L_1_out : std_logic := '0'; 
signal C_52_S_4_L_2_out : std_logic := '0'; 
signal C_52_S_4_L_3_out : std_logic := '0'; 
signal C_52_S_4_L_4_out : std_logic := '0'; 
signal C_52_S_4_L_5_out : std_logic := '0'; 
signal C_52_S_5_L_0_out : std_logic := '0'; 
signal C_52_S_5_L_1_out : std_logic := '0'; 
signal C_52_S_5_L_2_out : std_logic := '0'; 
signal C_52_S_5_L_3_out : std_logic := '0'; 
signal C_52_S_5_L_4_out : std_logic := '0'; 
signal C_52_S_5_L_5_out : std_logic := '0'; 
signal C_53_S_0_L_0_out : std_logic := '0'; 
signal C_53_S_0_L_1_out : std_logic := '0'; 
signal C_53_S_0_L_2_out : std_logic := '0'; 
signal C_53_S_0_L_3_out : std_logic := '0'; 
signal C_53_S_0_L_4_out : std_logic := '0'; 
signal C_53_S_0_L_5_out : std_logic := '0'; 
signal C_53_S_1_L_0_out : std_logic := '0'; 
signal C_53_S_1_L_1_out : std_logic := '0'; 
signal C_53_S_1_L_2_out : std_logic := '0'; 
signal C_53_S_1_L_3_out : std_logic := '0'; 
signal C_53_S_1_L_4_out : std_logic := '0'; 
signal C_53_S_1_L_5_out : std_logic := '0'; 
signal C_53_S_2_L_0_out : std_logic := '0'; 
signal C_53_S_2_L_1_out : std_logic := '0'; 
signal C_53_S_2_L_2_out : std_logic := '0'; 
signal C_53_S_2_L_3_out : std_logic := '0'; 
signal C_53_S_2_L_4_out : std_logic := '0'; 
signal C_53_S_2_L_5_out : std_logic := '0'; 
signal C_53_S_3_L_0_out : std_logic := '0'; 
signal C_53_S_3_L_1_out : std_logic := '0'; 
signal C_53_S_3_L_2_out : std_logic := '0'; 
signal C_53_S_3_L_3_out : std_logic := '0'; 
signal C_53_S_3_L_4_out : std_logic := '0'; 
signal C_53_S_3_L_5_out : std_logic := '0'; 
signal C_53_S_4_L_0_out : std_logic := '0'; 
signal C_53_S_4_L_1_out : std_logic := '0'; 
signal C_53_S_4_L_2_out : std_logic := '0'; 
signal C_53_S_4_L_3_out : std_logic := '0'; 
signal C_53_S_4_L_4_out : std_logic := '0'; 
signal C_53_S_4_L_5_out : std_logic := '0'; 
signal C_53_S_5_L_0_out : std_logic := '0'; 
signal C_53_S_5_L_1_out : std_logic := '0'; 
signal C_53_S_5_L_2_out : std_logic := '0'; 
signal C_53_S_5_L_3_out : std_logic := '0'; 
signal C_53_S_5_L_4_out : std_logic := '0'; 
signal C_53_S_5_L_5_out : std_logic := '0'; 
signal C_54_S_0_L_0_out : std_logic := '0'; 
signal C_54_S_0_L_1_out : std_logic := '0'; 
signal C_54_S_0_L_2_out : std_logic := '0'; 
signal C_54_S_0_L_3_out : std_logic := '0'; 
signal C_54_S_0_L_4_out : std_logic := '0'; 
signal C_54_S_0_L_5_out : std_logic := '0'; 
signal C_54_S_1_L_0_out : std_logic := '0'; 
signal C_54_S_1_L_1_out : std_logic := '0'; 
signal C_54_S_1_L_2_out : std_logic := '0'; 
signal C_54_S_1_L_3_out : std_logic := '0'; 
signal C_54_S_1_L_4_out : std_logic := '0'; 
signal C_54_S_1_L_5_out : std_logic := '0'; 
signal C_54_S_2_L_0_out : std_logic := '0'; 
signal C_54_S_2_L_1_out : std_logic := '0'; 
signal C_54_S_2_L_2_out : std_logic := '0'; 
signal C_54_S_2_L_3_out : std_logic := '0'; 
signal C_54_S_2_L_4_out : std_logic := '0'; 
signal C_54_S_2_L_5_out : std_logic := '0'; 
signal C_54_S_3_L_0_out : std_logic := '0'; 
signal C_54_S_3_L_1_out : std_logic := '0'; 
signal C_54_S_3_L_2_out : std_logic := '0'; 
signal C_54_S_3_L_3_out : std_logic := '0'; 
signal C_54_S_3_L_4_out : std_logic := '0'; 
signal C_54_S_3_L_5_out : std_logic := '0'; 
signal C_54_S_4_L_0_out : std_logic := '0'; 
signal C_54_S_4_L_1_out : std_logic := '0'; 
signal C_54_S_4_L_2_out : std_logic := '0'; 
signal C_54_S_4_L_3_out : std_logic := '0'; 
signal C_54_S_4_L_4_out : std_logic := '0'; 
signal C_54_S_4_L_5_out : std_logic := '0'; 
signal C_54_S_5_L_0_out : std_logic := '0'; 
signal C_54_S_5_L_1_out : std_logic := '0'; 
signal C_54_S_5_L_2_out : std_logic := '0'; 
signal C_54_S_5_L_3_out : std_logic := '0'; 
signal C_54_S_5_L_4_out : std_logic := '0'; 
signal C_54_S_5_L_5_out : std_logic := '0'; 
signal C_55_S_0_L_0_out : std_logic := '0'; 
signal C_55_S_0_L_1_out : std_logic := '0'; 
signal C_55_S_0_L_2_out : std_logic := '0'; 
signal C_55_S_0_L_3_out : std_logic := '0'; 
signal C_55_S_0_L_4_out : std_logic := '0'; 
signal C_55_S_0_L_5_out : std_logic := '0'; 
signal C_55_S_1_L_0_out : std_logic := '0'; 
signal C_55_S_1_L_1_out : std_logic := '0'; 
signal C_55_S_1_L_2_out : std_logic := '0'; 
signal C_55_S_1_L_3_out : std_logic := '0'; 
signal C_55_S_1_L_4_out : std_logic := '0'; 
signal C_55_S_1_L_5_out : std_logic := '0'; 
signal C_55_S_2_L_0_out : std_logic := '0'; 
signal C_55_S_2_L_1_out : std_logic := '0'; 
signal C_55_S_2_L_2_out : std_logic := '0'; 
signal C_55_S_2_L_3_out : std_logic := '0'; 
signal C_55_S_2_L_4_out : std_logic := '0'; 
signal C_55_S_2_L_5_out : std_logic := '0'; 
signal C_55_S_3_L_0_out : std_logic := '0'; 
signal C_55_S_3_L_1_out : std_logic := '0'; 
signal C_55_S_3_L_2_out : std_logic := '0'; 
signal C_55_S_3_L_3_out : std_logic := '0'; 
signal C_55_S_3_L_4_out : std_logic := '0'; 
signal C_55_S_3_L_5_out : std_logic := '0'; 
signal C_55_S_4_L_0_out : std_logic := '0'; 
signal C_55_S_4_L_1_out : std_logic := '0'; 
signal C_55_S_4_L_2_out : std_logic := '0'; 
signal C_55_S_4_L_3_out : std_logic := '0'; 
signal C_55_S_4_L_4_out : std_logic := '0'; 
signal C_55_S_4_L_5_out : std_logic := '0'; 
signal C_55_S_5_L_0_out : std_logic := '0'; 
signal C_55_S_5_L_1_out : std_logic := '0'; 
signal C_55_S_5_L_2_out : std_logic := '0'; 
signal C_55_S_5_L_3_out : std_logic := '0'; 
signal C_55_S_5_L_4_out : std_logic := '0'; 
signal C_55_S_5_L_5_out : std_logic := '0'; 
signal C_56_S_0_L_0_out : std_logic := '0'; 
signal C_56_S_0_L_1_out : std_logic := '0'; 
signal C_56_S_0_L_2_out : std_logic := '0'; 
signal C_56_S_0_L_3_out : std_logic := '0'; 
signal C_56_S_0_L_4_out : std_logic := '0'; 
signal C_56_S_0_L_5_out : std_logic := '0'; 
signal C_56_S_1_L_0_out : std_logic := '0'; 
signal C_56_S_1_L_1_out : std_logic := '0'; 
signal C_56_S_1_L_2_out : std_logic := '0'; 
signal C_56_S_1_L_3_out : std_logic := '0'; 
signal C_56_S_1_L_4_out : std_logic := '0'; 
signal C_56_S_1_L_5_out : std_logic := '0'; 
signal C_56_S_2_L_0_out : std_logic := '0'; 
signal C_56_S_2_L_1_out : std_logic := '0'; 
signal C_56_S_2_L_2_out : std_logic := '0'; 
signal C_56_S_2_L_3_out : std_logic := '0'; 
signal C_56_S_2_L_4_out : std_logic := '0'; 
signal C_56_S_2_L_5_out : std_logic := '0'; 
signal C_56_S_3_L_0_out : std_logic := '0'; 
signal C_56_S_3_L_1_out : std_logic := '0'; 
signal C_56_S_3_L_2_out : std_logic := '0'; 
signal C_56_S_3_L_3_out : std_logic := '0'; 
signal C_56_S_3_L_4_out : std_logic := '0'; 
signal C_56_S_3_L_5_out : std_logic := '0'; 
signal C_56_S_4_L_0_out : std_logic := '0'; 
signal C_56_S_4_L_1_out : std_logic := '0'; 
signal C_56_S_4_L_2_out : std_logic := '0'; 
signal C_56_S_4_L_3_out : std_logic := '0'; 
signal C_56_S_4_L_4_out : std_logic := '0'; 
signal C_56_S_4_L_5_out : std_logic := '0'; 
signal C_56_S_5_L_0_out : std_logic := '0'; 
signal C_56_S_5_L_1_out : std_logic := '0'; 
signal C_56_S_5_L_2_out : std_logic := '0'; 
signal C_56_S_5_L_3_out : std_logic := '0'; 
signal C_56_S_5_L_4_out : std_logic := '0'; 
signal C_56_S_5_L_5_out : std_logic := '0'; 
signal C_57_S_0_L_0_out : std_logic := '0'; 
signal C_57_S_0_L_1_out : std_logic := '0'; 
signal C_57_S_0_L_2_out : std_logic := '0'; 
signal C_57_S_0_L_3_out : std_logic := '0'; 
signal C_57_S_0_L_4_out : std_logic := '0'; 
signal C_57_S_0_L_5_out : std_logic := '0'; 
signal C_57_S_1_L_0_out : std_logic := '0'; 
signal C_57_S_1_L_1_out : std_logic := '0'; 
signal C_57_S_1_L_2_out : std_logic := '0'; 
signal C_57_S_1_L_3_out : std_logic := '0'; 
signal C_57_S_1_L_4_out : std_logic := '0'; 
signal C_57_S_1_L_5_out : std_logic := '0'; 
signal C_57_S_2_L_0_out : std_logic := '0'; 
signal C_57_S_2_L_1_out : std_logic := '0'; 
signal C_57_S_2_L_2_out : std_logic := '0'; 
signal C_57_S_2_L_3_out : std_logic := '0'; 
signal C_57_S_2_L_4_out : std_logic := '0'; 
signal C_57_S_2_L_5_out : std_logic := '0'; 
signal C_57_S_3_L_0_out : std_logic := '0'; 
signal C_57_S_3_L_1_out : std_logic := '0'; 
signal C_57_S_3_L_2_out : std_logic := '0'; 
signal C_57_S_3_L_3_out : std_logic := '0'; 
signal C_57_S_3_L_4_out : std_logic := '0'; 
signal C_57_S_3_L_5_out : std_logic := '0'; 
signal C_57_S_4_L_0_out : std_logic := '0'; 
signal C_57_S_4_L_1_out : std_logic := '0'; 
signal C_57_S_4_L_2_out : std_logic := '0'; 
signal C_57_S_4_L_3_out : std_logic := '0'; 
signal C_57_S_4_L_4_out : std_logic := '0'; 
signal C_57_S_4_L_5_out : std_logic := '0'; 
signal C_57_S_5_L_0_out : std_logic := '0'; 
signal C_57_S_5_L_1_out : std_logic := '0'; 
signal C_57_S_5_L_2_out : std_logic := '0'; 
signal C_57_S_5_L_3_out : std_logic := '0'; 
signal C_57_S_5_L_4_out : std_logic := '0'; 
signal C_57_S_5_L_5_out : std_logic := '0'; 
signal C_58_S_0_L_0_out : std_logic := '0'; 
signal C_58_S_0_L_1_out : std_logic := '0'; 
signal C_58_S_0_L_2_out : std_logic := '0'; 
signal C_58_S_0_L_3_out : std_logic := '0'; 
signal C_58_S_0_L_4_out : std_logic := '0'; 
signal C_58_S_0_L_5_out : std_logic := '0'; 
signal C_58_S_1_L_0_out : std_logic := '0'; 
signal C_58_S_1_L_1_out : std_logic := '0'; 
signal C_58_S_1_L_2_out : std_logic := '0'; 
signal C_58_S_1_L_3_out : std_logic := '0'; 
signal C_58_S_1_L_4_out : std_logic := '0'; 
signal C_58_S_1_L_5_out : std_logic := '0'; 
signal C_58_S_2_L_0_out : std_logic := '0'; 
signal C_58_S_2_L_1_out : std_logic := '0'; 
signal C_58_S_2_L_2_out : std_logic := '0'; 
signal C_58_S_2_L_3_out : std_logic := '0'; 
signal C_58_S_2_L_4_out : std_logic := '0'; 
signal C_58_S_2_L_5_out : std_logic := '0'; 
signal C_58_S_3_L_0_out : std_logic := '0'; 
signal C_58_S_3_L_1_out : std_logic := '0'; 
signal C_58_S_3_L_2_out : std_logic := '0'; 
signal C_58_S_3_L_3_out : std_logic := '0'; 
signal C_58_S_3_L_4_out : std_logic := '0'; 
signal C_58_S_3_L_5_out : std_logic := '0'; 
signal C_58_S_4_L_0_out : std_logic := '0'; 
signal C_58_S_4_L_1_out : std_logic := '0'; 
signal C_58_S_4_L_2_out : std_logic := '0'; 
signal C_58_S_4_L_3_out : std_logic := '0'; 
signal C_58_S_4_L_4_out : std_logic := '0'; 
signal C_58_S_4_L_5_out : std_logic := '0'; 
signal C_58_S_5_L_0_out : std_logic := '0'; 
signal C_58_S_5_L_1_out : std_logic := '0'; 
signal C_58_S_5_L_2_out : std_logic := '0'; 
signal C_58_S_5_L_3_out : std_logic := '0'; 
signal C_58_S_5_L_4_out : std_logic := '0'; 
signal C_58_S_5_L_5_out : std_logic := '0'; 
signal C_59_S_0_L_0_out : std_logic := '0'; 
signal C_59_S_0_L_1_out : std_logic := '0'; 
signal C_59_S_0_L_2_out : std_logic := '0'; 
signal C_59_S_0_L_3_out : std_logic := '0'; 
signal C_59_S_0_L_4_out : std_logic := '0'; 
signal C_59_S_0_L_5_out : std_logic := '0'; 
signal C_59_S_1_L_0_out : std_logic := '0'; 
signal C_59_S_1_L_1_out : std_logic := '0'; 
signal C_59_S_1_L_2_out : std_logic := '0'; 
signal C_59_S_1_L_3_out : std_logic := '0'; 
signal C_59_S_1_L_4_out : std_logic := '0'; 
signal C_59_S_1_L_5_out : std_logic := '0'; 
signal C_59_S_2_L_0_out : std_logic := '0'; 
signal C_59_S_2_L_1_out : std_logic := '0'; 
signal C_59_S_2_L_2_out : std_logic := '0'; 
signal C_59_S_2_L_3_out : std_logic := '0'; 
signal C_59_S_2_L_4_out : std_logic := '0'; 
signal C_59_S_2_L_5_out : std_logic := '0'; 
signal C_59_S_3_L_0_out : std_logic := '0'; 
signal C_59_S_3_L_1_out : std_logic := '0'; 
signal C_59_S_3_L_2_out : std_logic := '0'; 
signal C_59_S_3_L_3_out : std_logic := '0'; 
signal C_59_S_3_L_4_out : std_logic := '0'; 
signal C_59_S_3_L_5_out : std_logic := '0'; 
signal C_59_S_4_L_0_out : std_logic := '0'; 
signal C_59_S_4_L_1_out : std_logic := '0'; 
signal C_59_S_4_L_2_out : std_logic := '0'; 
signal C_59_S_4_L_3_out : std_logic := '0'; 
signal C_59_S_4_L_4_out : std_logic := '0'; 
signal C_59_S_4_L_5_out : std_logic := '0'; 
signal C_59_S_5_L_0_out : std_logic := '0'; 
signal C_59_S_5_L_1_out : std_logic := '0'; 
signal C_59_S_5_L_2_out : std_logic := '0'; 
signal C_59_S_5_L_3_out : std_logic := '0'; 
signal C_59_S_5_L_4_out : std_logic := '0'; 
signal C_59_S_5_L_5_out : std_logic := '0'; 

signal C_0_S_0_out : std_logic := '0'; 
signal C_0_S_1_out : std_logic := '0'; 
signal C_0_S_2_out : std_logic := '0'; 
signal C_0_S_3_out : std_logic := '0'; 
signal C_0_S_4_out : std_logic := '0'; 
signal C_0_S_5_out : std_logic := '0'; 
signal C_1_S_0_out : std_logic := '0'; 
signal C_1_S_1_out : std_logic := '0'; 
signal C_1_S_2_out : std_logic := '0'; 
signal C_1_S_3_out : std_logic := '0'; 
signal C_1_S_4_out : std_logic := '0'; 
signal C_1_S_5_out : std_logic := '0'; 
signal C_2_S_0_out : std_logic := '0'; 
signal C_2_S_1_out : std_logic := '0'; 
signal C_2_S_2_out : std_logic := '0'; 
signal C_2_S_3_out : std_logic := '0'; 
signal C_2_S_4_out : std_logic := '0'; 
signal C_2_S_5_out : std_logic := '0'; 
signal C_3_S_0_out : std_logic := '0'; 
signal C_3_S_1_out : std_logic := '0'; 
signal C_3_S_2_out : std_logic := '0'; 
signal C_3_S_3_out : std_logic := '0'; 
signal C_3_S_4_out : std_logic := '0'; 
signal C_3_S_5_out : std_logic := '0'; 
signal C_4_S_0_out : std_logic := '0'; 
signal C_4_S_1_out : std_logic := '0'; 
signal C_4_S_2_out : std_logic := '0'; 
signal C_4_S_3_out : std_logic := '0'; 
signal C_4_S_4_out : std_logic := '0'; 
signal C_4_S_5_out : std_logic := '0'; 
signal C_5_S_0_out : std_logic := '0'; 
signal C_5_S_1_out : std_logic := '0'; 
signal C_5_S_2_out : std_logic := '0'; 
signal C_5_S_3_out : std_logic := '0'; 
signal C_5_S_4_out : std_logic := '0'; 
signal C_5_S_5_out : std_logic := '0'; 
signal C_6_S_0_out : std_logic := '0'; 
signal C_6_S_1_out : std_logic := '0'; 
signal C_6_S_2_out : std_logic := '0'; 
signal C_6_S_3_out : std_logic := '0'; 
signal C_6_S_4_out : std_logic := '0'; 
signal C_6_S_5_out : std_logic := '0'; 
signal C_7_S_0_out : std_logic := '0'; 
signal C_7_S_1_out : std_logic := '0'; 
signal C_7_S_2_out : std_logic := '0'; 
signal C_7_S_3_out : std_logic := '0'; 
signal C_7_S_4_out : std_logic := '0'; 
signal C_7_S_5_out : std_logic := '0'; 
signal C_8_S_0_out : std_logic := '0'; 
signal C_8_S_1_out : std_logic := '0'; 
signal C_8_S_2_out : std_logic := '0'; 
signal C_8_S_3_out : std_logic := '0'; 
signal C_8_S_4_out : std_logic := '0'; 
signal C_8_S_5_out : std_logic := '0'; 
signal C_9_S_0_out : std_logic := '0'; 
signal C_9_S_1_out : std_logic := '0'; 
signal C_9_S_2_out : std_logic := '0'; 
signal C_9_S_3_out : std_logic := '0'; 
signal C_9_S_4_out : std_logic := '0'; 
signal C_9_S_5_out : std_logic := '0'; 
signal C_10_S_0_out : std_logic := '0'; 
signal C_10_S_1_out : std_logic := '0'; 
signal C_10_S_2_out : std_logic := '0'; 
signal C_10_S_3_out : std_logic := '0'; 
signal C_10_S_4_out : std_logic := '0'; 
signal C_10_S_5_out : std_logic := '0'; 
signal C_11_S_0_out : std_logic := '0'; 
signal C_11_S_1_out : std_logic := '0'; 
signal C_11_S_2_out : std_logic := '0'; 
signal C_11_S_3_out : std_logic := '0'; 
signal C_11_S_4_out : std_logic := '0'; 
signal C_11_S_5_out : std_logic := '0'; 
signal C_12_S_0_out : std_logic := '0'; 
signal C_12_S_1_out : std_logic := '0'; 
signal C_12_S_2_out : std_logic := '0'; 
signal C_12_S_3_out : std_logic := '0'; 
signal C_12_S_4_out : std_logic := '0'; 
signal C_12_S_5_out : std_logic := '0'; 
signal C_13_S_0_out : std_logic := '0'; 
signal C_13_S_1_out : std_logic := '0'; 
signal C_13_S_2_out : std_logic := '0'; 
signal C_13_S_3_out : std_logic := '0'; 
signal C_13_S_4_out : std_logic := '0'; 
signal C_13_S_5_out : std_logic := '0'; 
signal C_14_S_0_out : std_logic := '0'; 
signal C_14_S_1_out : std_logic := '0'; 
signal C_14_S_2_out : std_logic := '0'; 
signal C_14_S_3_out : std_logic := '0'; 
signal C_14_S_4_out : std_logic := '0'; 
signal C_14_S_5_out : std_logic := '0'; 
signal C_15_S_0_out : std_logic := '0'; 
signal C_15_S_1_out : std_logic := '0'; 
signal C_15_S_2_out : std_logic := '0'; 
signal C_15_S_3_out : std_logic := '0'; 
signal C_15_S_4_out : std_logic := '0'; 
signal C_15_S_5_out : std_logic := '0'; 
signal C_16_S_0_out : std_logic := '0'; 
signal C_16_S_1_out : std_logic := '0'; 
signal C_16_S_2_out : std_logic := '0'; 
signal C_16_S_3_out : std_logic := '0'; 
signal C_16_S_4_out : std_logic := '0'; 
signal C_16_S_5_out : std_logic := '0'; 
signal C_17_S_0_out : std_logic := '0'; 
signal C_17_S_1_out : std_logic := '0'; 
signal C_17_S_2_out : std_logic := '0'; 
signal C_17_S_3_out : std_logic := '0'; 
signal C_17_S_4_out : std_logic := '0'; 
signal C_17_S_5_out : std_logic := '0'; 
signal C_18_S_0_out : std_logic := '0'; 
signal C_18_S_1_out : std_logic := '0'; 
signal C_18_S_2_out : std_logic := '0'; 
signal C_18_S_3_out : std_logic := '0'; 
signal C_18_S_4_out : std_logic := '0'; 
signal C_18_S_5_out : std_logic := '0'; 
signal C_19_S_0_out : std_logic := '0'; 
signal C_19_S_1_out : std_logic := '0'; 
signal C_19_S_2_out : std_logic := '0'; 
signal C_19_S_3_out : std_logic := '0'; 
signal C_19_S_4_out : std_logic := '0'; 
signal C_19_S_5_out : std_logic := '0'; 
signal C_20_S_0_out : std_logic := '0'; 
signal C_20_S_1_out : std_logic := '0'; 
signal C_20_S_2_out : std_logic := '0'; 
signal C_20_S_3_out : std_logic := '0'; 
signal C_20_S_4_out : std_logic := '0'; 
signal C_20_S_5_out : std_logic := '0'; 
signal C_21_S_0_out : std_logic := '0'; 
signal C_21_S_1_out : std_logic := '0'; 
signal C_21_S_2_out : std_logic := '0'; 
signal C_21_S_3_out : std_logic := '0'; 
signal C_21_S_4_out : std_logic := '0'; 
signal C_21_S_5_out : std_logic := '0'; 
signal C_22_S_0_out : std_logic := '0'; 
signal C_22_S_1_out : std_logic := '0'; 
signal C_22_S_2_out : std_logic := '0'; 
signal C_22_S_3_out : std_logic := '0'; 
signal C_22_S_4_out : std_logic := '0'; 
signal C_22_S_5_out : std_logic := '0'; 
signal C_23_S_0_out : std_logic := '0'; 
signal C_23_S_1_out : std_logic := '0'; 
signal C_23_S_2_out : std_logic := '0'; 
signal C_23_S_3_out : std_logic := '0'; 
signal C_23_S_4_out : std_logic := '0'; 
signal C_23_S_5_out : std_logic := '0'; 
signal C_24_S_0_out : std_logic := '0'; 
signal C_24_S_1_out : std_logic := '0'; 
signal C_24_S_2_out : std_logic := '0'; 
signal C_24_S_3_out : std_logic := '0'; 
signal C_24_S_4_out : std_logic := '0'; 
signal C_24_S_5_out : std_logic := '0'; 
signal C_25_S_0_out : std_logic := '0'; 
signal C_25_S_1_out : std_logic := '0'; 
signal C_25_S_2_out : std_logic := '0'; 
signal C_25_S_3_out : std_logic := '0'; 
signal C_25_S_4_out : std_logic := '0'; 
signal C_25_S_5_out : std_logic := '0'; 
signal C_26_S_0_out : std_logic := '0'; 
signal C_26_S_1_out : std_logic := '0'; 
signal C_26_S_2_out : std_logic := '0'; 
signal C_26_S_3_out : std_logic := '0'; 
signal C_26_S_4_out : std_logic := '0'; 
signal C_26_S_5_out : std_logic := '0'; 
signal C_27_S_0_out : std_logic := '0'; 
signal C_27_S_1_out : std_logic := '0'; 
signal C_27_S_2_out : std_logic := '0'; 
signal C_27_S_3_out : std_logic := '0'; 
signal C_27_S_4_out : std_logic := '0'; 
signal C_27_S_5_out : std_logic := '0'; 
signal C_28_S_0_out : std_logic := '0'; 
signal C_28_S_1_out : std_logic := '0'; 
signal C_28_S_2_out : std_logic := '0'; 
signal C_28_S_3_out : std_logic := '0'; 
signal C_28_S_4_out : std_logic := '0'; 
signal C_28_S_5_out : std_logic := '0'; 
signal C_29_S_0_out : std_logic := '0'; 
signal C_29_S_1_out : std_logic := '0'; 
signal C_29_S_2_out : std_logic := '0'; 
signal C_29_S_3_out : std_logic := '0'; 
signal C_29_S_4_out : std_logic := '0'; 
signal C_29_S_5_out : std_logic := '0'; 
signal C_30_S_0_out : std_logic := '0'; 
signal C_30_S_1_out : std_logic := '0'; 
signal C_30_S_2_out : std_logic := '0'; 
signal C_30_S_3_out : std_logic := '0'; 
signal C_30_S_4_out : std_logic := '0'; 
signal C_30_S_5_out : std_logic := '0'; 
signal C_31_S_0_out : std_logic := '0'; 
signal C_31_S_1_out : std_logic := '0'; 
signal C_31_S_2_out : std_logic := '0'; 
signal C_31_S_3_out : std_logic := '0'; 
signal C_31_S_4_out : std_logic := '0'; 
signal C_31_S_5_out : std_logic := '0'; 
signal C_32_S_0_out : std_logic := '0'; 
signal C_32_S_1_out : std_logic := '0'; 
signal C_32_S_2_out : std_logic := '0'; 
signal C_32_S_3_out : std_logic := '0'; 
signal C_32_S_4_out : std_logic := '0'; 
signal C_32_S_5_out : std_logic := '0'; 
signal C_33_S_0_out : std_logic := '0'; 
signal C_33_S_1_out : std_logic := '0'; 
signal C_33_S_2_out : std_logic := '0'; 
signal C_33_S_3_out : std_logic := '0'; 
signal C_33_S_4_out : std_logic := '0'; 
signal C_33_S_5_out : std_logic := '0'; 
signal C_34_S_0_out : std_logic := '0'; 
signal C_34_S_1_out : std_logic := '0'; 
signal C_34_S_2_out : std_logic := '0'; 
signal C_34_S_3_out : std_logic := '0'; 
signal C_34_S_4_out : std_logic := '0'; 
signal C_34_S_5_out : std_logic := '0'; 
signal C_35_S_0_out : std_logic := '0'; 
signal C_35_S_1_out : std_logic := '0'; 
signal C_35_S_2_out : std_logic := '0'; 
signal C_35_S_3_out : std_logic := '0'; 
signal C_35_S_4_out : std_logic := '0'; 
signal C_35_S_5_out : std_logic := '0'; 
signal C_36_S_0_out : std_logic := '0'; 
signal C_36_S_1_out : std_logic := '0'; 
signal C_36_S_2_out : std_logic := '0'; 
signal C_36_S_3_out : std_logic := '0'; 
signal C_36_S_4_out : std_logic := '0'; 
signal C_36_S_5_out : std_logic := '0'; 
signal C_37_S_0_out : std_logic := '0'; 
signal C_37_S_1_out : std_logic := '0'; 
signal C_37_S_2_out : std_logic := '0'; 
signal C_37_S_3_out : std_logic := '0'; 
signal C_37_S_4_out : std_logic := '0'; 
signal C_37_S_5_out : std_logic := '0'; 
signal C_38_S_0_out : std_logic := '0'; 
signal C_38_S_1_out : std_logic := '0'; 
signal C_38_S_2_out : std_logic := '0'; 
signal C_38_S_3_out : std_logic := '0'; 
signal C_38_S_4_out : std_logic := '0'; 
signal C_38_S_5_out : std_logic := '0'; 
signal C_39_S_0_out : std_logic := '0'; 
signal C_39_S_1_out : std_logic := '0'; 
signal C_39_S_2_out : std_logic := '0'; 
signal C_39_S_3_out : std_logic := '0'; 
signal C_39_S_4_out : std_logic := '0'; 
signal C_39_S_5_out : std_logic := '0'; 
signal C_40_S_0_out : std_logic := '0'; 
signal C_40_S_1_out : std_logic := '0'; 
signal C_40_S_2_out : std_logic := '0'; 
signal C_40_S_3_out : std_logic := '0'; 
signal C_40_S_4_out : std_logic := '0'; 
signal C_40_S_5_out : std_logic := '0'; 
signal C_41_S_0_out : std_logic := '0'; 
signal C_41_S_1_out : std_logic := '0'; 
signal C_41_S_2_out : std_logic := '0'; 
signal C_41_S_3_out : std_logic := '0'; 
signal C_41_S_4_out : std_logic := '0'; 
signal C_41_S_5_out : std_logic := '0'; 
signal C_42_S_0_out : std_logic := '0'; 
signal C_42_S_1_out : std_logic := '0'; 
signal C_42_S_2_out : std_logic := '0'; 
signal C_42_S_3_out : std_logic := '0'; 
signal C_42_S_4_out : std_logic := '0'; 
signal C_42_S_5_out : std_logic := '0'; 
signal C_43_S_0_out : std_logic := '0'; 
signal C_43_S_1_out : std_logic := '0'; 
signal C_43_S_2_out : std_logic := '0'; 
signal C_43_S_3_out : std_logic := '0'; 
signal C_43_S_4_out : std_logic := '0'; 
signal C_43_S_5_out : std_logic := '0'; 
signal C_44_S_0_out : std_logic := '0'; 
signal C_44_S_1_out : std_logic := '0'; 
signal C_44_S_2_out : std_logic := '0'; 
signal C_44_S_3_out : std_logic := '0'; 
signal C_44_S_4_out : std_logic := '0'; 
signal C_44_S_5_out : std_logic := '0'; 
signal C_45_S_0_out : std_logic := '0'; 
signal C_45_S_1_out : std_logic := '0'; 
signal C_45_S_2_out : std_logic := '0'; 
signal C_45_S_3_out : std_logic := '0'; 
signal C_45_S_4_out : std_logic := '0'; 
signal C_45_S_5_out : std_logic := '0'; 
signal C_46_S_0_out : std_logic := '0'; 
signal C_46_S_1_out : std_logic := '0'; 
signal C_46_S_2_out : std_logic := '0'; 
signal C_46_S_3_out : std_logic := '0'; 
signal C_46_S_4_out : std_logic := '0'; 
signal C_46_S_5_out : std_logic := '0'; 
signal C_47_S_0_out : std_logic := '0'; 
signal C_47_S_1_out : std_logic := '0'; 
signal C_47_S_2_out : std_logic := '0'; 
signal C_47_S_3_out : std_logic := '0'; 
signal C_47_S_4_out : std_logic := '0'; 
signal C_47_S_5_out : std_logic := '0'; 
signal C_48_S_0_out : std_logic := '0'; 
signal C_48_S_1_out : std_logic := '0'; 
signal C_48_S_2_out : std_logic := '0'; 
signal C_48_S_3_out : std_logic := '0'; 
signal C_48_S_4_out : std_logic := '0'; 
signal C_48_S_5_out : std_logic := '0'; 
signal C_49_S_0_out : std_logic := '0'; 
signal C_49_S_1_out : std_logic := '0'; 
signal C_49_S_2_out : std_logic := '0'; 
signal C_49_S_3_out : std_logic := '0'; 
signal C_49_S_4_out : std_logic := '0'; 
signal C_49_S_5_out : std_logic := '0'; 
signal C_50_S_0_out : std_logic := '0'; 
signal C_50_S_1_out : std_logic := '0'; 
signal C_50_S_2_out : std_logic := '0'; 
signal C_50_S_3_out : std_logic := '0'; 
signal C_50_S_4_out : std_logic := '0'; 
signal C_50_S_5_out : std_logic := '0'; 
signal C_51_S_0_out : std_logic := '0'; 
signal C_51_S_1_out : std_logic := '0'; 
signal C_51_S_2_out : std_logic := '0'; 
signal C_51_S_3_out : std_logic := '0'; 
signal C_51_S_4_out : std_logic := '0'; 
signal C_51_S_5_out : std_logic := '0'; 
signal C_52_S_0_out : std_logic := '0'; 
signal C_52_S_1_out : std_logic := '0'; 
signal C_52_S_2_out : std_logic := '0'; 
signal C_52_S_3_out : std_logic := '0'; 
signal C_52_S_4_out : std_logic := '0'; 
signal C_52_S_5_out : std_logic := '0'; 
signal C_53_S_0_out : std_logic := '0'; 
signal C_53_S_1_out : std_logic := '0'; 
signal C_53_S_2_out : std_logic := '0'; 
signal C_53_S_3_out : std_logic := '0'; 
signal C_53_S_4_out : std_logic := '0'; 
signal C_53_S_5_out : std_logic := '0'; 
signal C_54_S_0_out : std_logic := '0'; 
signal C_54_S_1_out : std_logic := '0'; 
signal C_54_S_2_out : std_logic := '0'; 
signal C_54_S_3_out : std_logic := '0'; 
signal C_54_S_4_out : std_logic := '0'; 
signal C_54_S_5_out : std_logic := '0'; 
signal C_55_S_0_out : std_logic := '0'; 
signal C_55_S_1_out : std_logic := '0'; 
signal C_55_S_2_out : std_logic := '0'; 
signal C_55_S_3_out : std_logic := '0'; 
signal C_55_S_4_out : std_logic := '0'; 
signal C_55_S_5_out : std_logic := '0'; 
signal C_56_S_0_out : std_logic := '0'; 
signal C_56_S_1_out : std_logic := '0'; 
signal C_56_S_2_out : std_logic := '0'; 
signal C_56_S_3_out : std_logic := '0'; 
signal C_56_S_4_out : std_logic := '0'; 
signal C_56_S_5_out : std_logic := '0'; 
signal C_57_S_0_out : std_logic := '0'; 
signal C_57_S_1_out : std_logic := '0'; 
signal C_57_S_2_out : std_logic := '0'; 
signal C_57_S_3_out : std_logic := '0'; 
signal C_57_S_4_out : std_logic := '0'; 
signal C_57_S_5_out : std_logic := '0'; 
signal C_58_S_0_out : std_logic := '0'; 
signal C_58_S_1_out : std_logic := '0'; 
signal C_58_S_2_out : std_logic := '0'; 
signal C_58_S_3_out : std_logic := '0'; 
signal C_58_S_4_out : std_logic := '0'; 
signal C_58_S_5_out : std_logic := '0'; 
signal C_59_S_0_out : std_logic := '0'; 
signal C_59_S_1_out : std_logic := '0'; 
signal C_59_S_2_out : std_logic := '0'; 
signal C_59_S_3_out : std_logic := '0'; 
signal C_59_S_4_out : std_logic := '0'; 
signal C_59_S_5_out : std_logic := '0'; signal C_0_B_7_out : std_logic := '0'; 
 signal C_0_B_6_out : std_logic := '0'; 
 signal C_0_B_5_out : std_logic := '0'; 
 signal C_0_B_4_out : std_logic := '0'; 
 signal C_0_B_3_out : std_logic := '0'; 
 signal C_0_B_2_out : std_logic := '0'; 
 signal C_0_B_1_out : std_logic := '0'; 
 signal C_0_B_0_out : std_logic := '0'; 
 signal C_1_B_7_out : std_logic := '0'; 
 signal C_1_B_6_out : std_logic := '0'; 
 signal C_1_B_5_out : std_logic := '0'; 
 signal C_1_B_4_out : std_logic := '0'; 
 signal C_1_B_3_out : std_logic := '0'; 
 signal C_1_B_2_out : std_logic := '0'; 
 signal C_1_B_1_out : std_logic := '0'; 
 signal C_1_B_0_out : std_logic := '0'; 
 signal C_2_B_7_out : std_logic := '0'; 
 signal C_2_B_6_out : std_logic := '0'; 
 signal C_2_B_5_out : std_logic := '0'; 
 signal C_2_B_4_out : std_logic := '0'; 
 signal C_2_B_3_out : std_logic := '0'; 
 signal C_2_B_2_out : std_logic := '0'; 
 signal C_2_B_1_out : std_logic := '0'; 
 signal C_2_B_0_out : std_logic := '0'; 
 signal C_3_B_7_out : std_logic := '0'; 
 signal C_3_B_6_out : std_logic := '0'; 
 signal C_3_B_5_out : std_logic := '0'; 
 signal C_3_B_4_out : std_logic := '0'; 
 signal C_3_B_3_out : std_logic := '0'; 
 signal C_3_B_2_out : std_logic := '0'; 
 signal C_3_B_1_out : std_logic := '0'; 
 signal C_3_B_0_out : std_logic := '0'; 
 signal C_4_B_7_out : std_logic := '0'; 
 signal C_4_B_6_out : std_logic := '0'; 
 signal C_4_B_5_out : std_logic := '0'; 
 signal C_4_B_4_out : std_logic := '0'; 
 signal C_4_B_3_out : std_logic := '0'; 
 signal C_4_B_2_out : std_logic := '0'; 
 signal C_4_B_1_out : std_logic := '0'; 
 signal C_4_B_0_out : std_logic := '0'; 
 signal C_5_B_7_out : std_logic := '0'; 
 signal C_5_B_6_out : std_logic := '0'; 
 signal C_5_B_5_out : std_logic := '0'; 
 signal C_5_B_4_out : std_logic := '0'; 
 signal C_5_B_3_out : std_logic := '0'; 
 signal C_5_B_2_out : std_logic := '0'; 
 signal C_5_B_1_out : std_logic := '0'; 
 signal C_5_B_0_out : std_logic := '0'; 
 signal C_6_B_7_out : std_logic := '0'; 
 signal C_6_B_6_out : std_logic := '0'; 
 signal C_6_B_5_out : std_logic := '0'; 
 signal C_6_B_4_out : std_logic := '0'; 
 signal C_6_B_3_out : std_logic := '0'; 
 signal C_6_B_2_out : std_logic := '0'; 
 signal C_6_B_1_out : std_logic := '0'; 
 signal C_6_B_0_out : std_logic := '0'; 
 signal C_7_B_7_out : std_logic := '0'; 
 signal C_7_B_6_out : std_logic := '0'; 
 signal C_7_B_5_out : std_logic := '0'; 
 signal C_7_B_4_out : std_logic := '0'; 
 signal C_7_B_3_out : std_logic := '0'; 
 signal C_7_B_2_out : std_logic := '0'; 
 signal C_7_B_1_out : std_logic := '0'; 
 signal C_7_B_0_out : std_logic := '0'; 
 signal C_8_B_7_out : std_logic := '0'; 
 signal C_8_B_6_out : std_logic := '0'; 
 signal C_8_B_5_out : std_logic := '0'; 
 signal C_8_B_4_out : std_logic := '0'; 
 signal C_8_B_3_out : std_logic := '0'; 
 signal C_8_B_2_out : std_logic := '0'; 
 signal C_8_B_1_out : std_logic := '0'; 
 signal C_8_B_0_out : std_logic := '0'; 
 signal C_9_B_7_out : std_logic := '0'; 
 signal C_9_B_6_out : std_logic := '0'; 
 signal C_9_B_5_out : std_logic := '0'; 
 signal C_9_B_4_out : std_logic := '0'; 
 signal C_9_B_3_out : std_logic := '0'; 
 signal C_9_B_2_out : std_logic := '0'; 
 signal C_9_B_1_out : std_logic := '0'; 
 signal C_9_B_0_out : std_logic := '0'; 


begin


C_0_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111101110111111111000000011111110111110001111000000000000") port map( O =>C_0_S_0_L_0_out, I0 =>  inp_feat(234), I1 =>  inp_feat(435), I2 =>  inp_feat(82), I3 =>  inp_feat(0), I4 =>  inp_feat(102), I5 =>  inp_feat(327)); 
C_0_S_0_L_1_inst : LUT6 generic map(INIT => "1111001011010011000000000101010111110111111000101100111111111101") port map( O =>C_0_S_0_L_1_out, I0 =>  inp_feat(173), I1 =>  inp_feat(160), I2 =>  inp_feat(71), I3 =>  inp_feat(323), I4 =>  inp_feat(497), I5 =>  inp_feat(419)); 
C_0_S_0_L_2_inst : LUT6 generic map(INIT => "0101000101010100001010101011110011111001111101000110100011111100") port map( O =>C_0_S_0_L_2_out, I0 =>  inp_feat(27), I1 =>  inp_feat(153), I2 =>  inp_feat(15), I3 =>  inp_feat(348), I4 =>  inp_feat(392), I5 =>  inp_feat(419)); 
C_0_S_0_L_3_inst : LUT6 generic map(INIT => "1111111111101110101101110010111001101011000011010011010110100000") port map( O =>C_0_S_0_L_3_out, I0 =>  inp_feat(420), I1 =>  inp_feat(373), I2 =>  inp_feat(71), I3 =>  inp_feat(151), I4 =>  inp_feat(74), I5 =>  inp_feat(82)); 
C_0_S_0_L_4_inst : LUT6 generic map(INIT => "0100011000000011111011100000011111110011111000111111111111110000") port map( O =>C_0_S_0_L_4_out, I0 =>  inp_feat(155), I1 =>  inp_feat(39), I2 =>  inp_feat(370), I3 =>  inp_feat(404), I4 =>  inp_feat(89), I5 =>  inp_feat(125)); 
C_0_S_0_L_5_inst : LUT6 generic map(INIT => "1111101011110010101111011110111011111011111111101111111001111111") port map( O =>C_0_S_0_L_5_out, I0 =>  inp_feat(338), I1 =>  inp_feat(133), I2 =>  inp_feat(50), I3 =>  inp_feat(404), I4 =>  inp_feat(309), I5 =>  inp_feat(16)); 
C_0_S_1_L_0_inst : LUT6 generic map(INIT => "1111001011010011000000000101010111110111111000101100111111111101") port map( O =>C_0_S_1_L_0_out, I0 =>  inp_feat(173), I1 =>  inp_feat(160), I2 =>  inp_feat(71), I3 =>  inp_feat(323), I4 =>  inp_feat(497), I5 =>  inp_feat(419)); 
C_0_S_1_L_1_inst : LUT6 generic map(INIT => "0101000101010100001010101011110011111001111101000110100011111100") port map( O =>C_0_S_1_L_1_out, I0 =>  inp_feat(27), I1 =>  inp_feat(153), I2 =>  inp_feat(15), I3 =>  inp_feat(348), I4 =>  inp_feat(392), I5 =>  inp_feat(419)); 
C_0_S_1_L_2_inst : LUT6 generic map(INIT => "1111111111101110101101110010111001101011000011010011010110100000") port map( O =>C_0_S_1_L_2_out, I0 =>  inp_feat(420), I1 =>  inp_feat(373), I2 =>  inp_feat(71), I3 =>  inp_feat(151), I4 =>  inp_feat(74), I5 =>  inp_feat(82)); 
C_0_S_1_L_3_inst : LUT6 generic map(INIT => "0100011000000011111011100000011111110011111000111111111111110000") port map( O =>C_0_S_1_L_3_out, I0 =>  inp_feat(155), I1 =>  inp_feat(39), I2 =>  inp_feat(370), I3 =>  inp_feat(404), I4 =>  inp_feat(89), I5 =>  inp_feat(125)); 
C_0_S_1_L_4_inst : LUT6 generic map(INIT => "1111101011110010101111011110111011111011111111101111111001111111") port map( O =>C_0_S_1_L_4_out, I0 =>  inp_feat(338), I1 =>  inp_feat(133), I2 =>  inp_feat(50), I3 =>  inp_feat(404), I4 =>  inp_feat(309), I5 =>  inp_feat(16)); 
C_0_S_1_L_5_inst : LUT6 generic map(INIT => "0001011000100001111111010100110111111111111010101111111101111111") port map( O =>C_0_S_1_L_5_out, I0 =>  inp_feat(155), I1 =>  inp_feat(133), I2 =>  inp_feat(50), I3 =>  inp_feat(404), I4 =>  inp_feat(309), I5 =>  inp_feat(16)); 
C_0_S_2_L_0_inst : LUT6 generic map(INIT => "0000101100110111000010111111101111110110111110000011010011111100") port map( O =>C_0_S_2_L_0_out, I0 =>  inp_feat(105), I1 =>  inp_feat(352), I2 =>  inp_feat(501), I3 =>  inp_feat(11), I4 =>  inp_feat(391), I5 =>  inp_feat(169)); 
C_0_S_2_L_1_inst : LUT6 generic map(INIT => "1101111000001110110111000000100011111111100110011110100010001000") port map( O =>C_0_S_2_L_1_out, I0 =>  inp_feat(418), I1 =>  inp_feat(74), I2 =>  inp_feat(10), I3 =>  inp_feat(488), I4 =>  inp_feat(208), I5 =>  inp_feat(507)); 
C_0_S_2_L_2_inst : LUT6 generic map(INIT => "0111000100110100000000100001111011111111101111101110111011101010") port map( O =>C_0_S_2_L_2_out, I0 =>  inp_feat(432), I1 =>  inp_feat(429), I2 =>  inp_feat(234), I3 =>  inp_feat(378), I4 =>  inp_feat(208), I5 =>  inp_feat(507)); 
C_0_S_2_L_3_inst : LUT6 generic map(INIT => "1101100000011011001011001100110011111001111101101111111010001010") port map( O =>C_0_S_2_L_3_out, I0 =>  inp_feat(458), I1 =>  inp_feat(350), I2 =>  inp_feat(169), I3 =>  inp_feat(156), I4 =>  inp_feat(211), I5 =>  inp_feat(175)); 
C_0_S_2_L_4_inst : LUT6 generic map(INIT => "0001111100010111010010010101110110111111010101111111111001011111") port map( O =>C_0_S_2_L_4_out, I0 =>  inp_feat(168), I1 =>  inp_feat(480), I2 =>  inp_feat(306), I3 =>  inp_feat(439), I4 =>  inp_feat(323), I5 =>  inp_feat(417)); 
C_0_S_2_L_5_inst : LUT6 generic map(INIT => "1100010110001000110011100010111111011111111101111111111100111010") port map( O =>C_0_S_2_L_5_out, I0 =>  inp_feat(389), I1 =>  inp_feat(467), I2 =>  inp_feat(29), I3 =>  inp_feat(34), I4 =>  inp_feat(89), I5 =>  inp_feat(125)); 
C_0_S_3_L_0_inst : LUT6 generic map(INIT => "1110111011110101111111101111101001001100011011110111001000000000") port map( O =>C_0_S_3_L_0_out, I0 =>  inp_feat(86), I1 =>  inp_feat(510), I2 =>  inp_feat(419), I3 =>  inp_feat(128), I4 =>  inp_feat(29), I5 =>  inp_feat(58)); 
C_0_S_3_L_1_inst : LUT6 generic map(INIT => "0100001000001100011110101011100011111101111101111110111111001000") port map( O =>C_0_S_3_L_1_out, I0 =>  inp_feat(106), I1 =>  inp_feat(95), I2 =>  inp_feat(501), I3 =>  inp_feat(313), I4 =>  inp_feat(211), I5 =>  inp_feat(175)); 
C_0_S_3_L_2_inst : LUT6 generic map(INIT => "0101011101110011110000110111000111111111111000101101110111100000") port map( O =>C_0_S_3_L_2_out, I0 =>  inp_feat(446), I1 =>  inp_feat(306), I2 =>  inp_feat(130), I3 =>  inp_feat(171), I4 =>  inp_feat(370), I5 =>  inp_feat(70)); 
C_0_S_3_L_3_inst : LUT6 generic map(INIT => "1100011110001110110100010001110110101111111111111101111111111111") port map( O =>C_0_S_3_L_3_out, I0 =>  inp_feat(373), I1 =>  inp_feat(2), I2 =>  inp_feat(77), I3 =>  inp_feat(363), I4 =>  inp_feat(476), I5 =>  inp_feat(66)); 
C_0_S_3_L_4_inst : LUT6 generic map(INIT => "1111011011111110101111111111000000000000111100001111111101110000") port map( O =>C_0_S_3_L_4_out, I0 =>  inp_feat(145), I1 =>  inp_feat(89), I2 =>  inp_feat(164), I3 =>  inp_feat(220), I4 =>  inp_feat(125), I5 =>  inp_feat(480)); 
C_0_S_3_L_5_inst : LUT6 generic map(INIT => "0011001001001110010111101110111100000110000011100000110111010111") port map( O =>C_0_S_3_L_5_out, I0 =>  inp_feat(11), I1 =>  inp_feat(77), I2 =>  inp_feat(174), I3 =>  inp_feat(417), I4 =>  inp_feat(94), I5 =>  inp_feat(25)); 
C_0_S_4_L_0_inst : LUT6 generic map(INIT => "1111110011101000101011001100000011111110111010111111110011110000") port map( O =>C_0_S_4_L_0_out, I0 =>  inp_feat(348), I1 =>  inp_feat(170), I2 =>  inp_feat(159), I3 =>  inp_feat(325), I4 =>  inp_feat(490), I5 =>  inp_feat(139)); 
C_0_S_4_L_1_inst : LUT6 generic map(INIT => "0000010000111011000011100011110110101111111011111011110111111111") port map( O =>C_0_S_4_L_1_out, I0 =>  inp_feat(346), I1 =>  inp_feat(102), I2 =>  inp_feat(375), I3 =>  inp_feat(363), I4 =>  inp_feat(476), I5 =>  inp_feat(66)); 
C_0_S_4_L_2_inst : LUT6 generic map(INIT => "1100110111111110100101101111101000001101010111010100000011110000") port map( O =>C_0_S_4_L_2_out, I0 =>  inp_feat(167), I1 =>  inp_feat(451), I2 =>  inp_feat(148), I3 =>  inp_feat(372), I4 =>  inp_feat(464), I5 =>  inp_feat(436)); 
C_0_S_4_L_3_inst : LUT6 generic map(INIT => "1110001010110010111001101010111101001100111110000100110011111110") port map( O =>C_0_S_4_L_3_out, I0 =>  inp_feat(435), I1 =>  inp_feat(31), I2 =>  inp_feat(234), I3 =>  inp_feat(327), I4 =>  inp_feat(373), I5 =>  inp_feat(445)); 
C_0_S_4_L_4_inst : LUT6 generic map(INIT => "0100110001111111000011110101110111101110111010000010010010101010") port map( O =>C_0_S_4_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(283), I2 =>  inp_feat(10), I3 =>  inp_feat(415), I4 =>  inp_feat(78), I5 =>  inp_feat(453)); 
C_0_S_4_L_5_inst : LUT6 generic map(INIT => "1111111101111111011001111110111100010111001011110111111111111111") port map( O =>C_0_S_4_L_5_out, I0 =>  inp_feat(510), I1 =>  inp_feat(262), I2 =>  inp_feat(383), I3 =>  inp_feat(274), I4 =>  inp_feat(484), I5 =>  inp_feat(105)); 
C_0_S_5_L_0_inst : LUT6 generic map(INIT => "0000010000111001000011100011110110101111111011111011110111111111") port map( O =>C_0_S_5_L_0_out, I0 =>  inp_feat(346), I1 =>  inp_feat(102), I2 =>  inp_feat(375), I3 =>  inp_feat(363), I4 =>  inp_feat(476), I5 =>  inp_feat(66)); 
C_0_S_5_L_1_inst : LUT6 generic map(INIT => "1111001110001111111011011000111110111011101011011111111111101111") port map( O =>C_0_S_5_L_1_out, I0 =>  inp_feat(160), I1 =>  inp_feat(446), I2 =>  inp_feat(29), I3 =>  inp_feat(114), I4 =>  inp_feat(89), I5 =>  inp_feat(125)); 
C_0_S_5_L_2_inst : LUT6 generic map(INIT => "0100010111010001110100111101010111111101111101101111110101111101") port map( O =>C_0_S_5_L_2_out, I0 =>  inp_feat(29), I1 =>  inp_feat(432), I2 =>  inp_feat(250), I3 =>  inp_feat(178), I4 =>  inp_feat(89), I5 =>  inp_feat(125)); 
C_0_S_5_L_3_inst : LUT6 generic map(INIT => "0010110010101000111111001100110011101101110011111110111111111111") port map( O =>C_0_S_5_L_3_out, I0 =>  inp_feat(403), I1 =>  inp_feat(370), I2 =>  inp_feat(174), I3 =>  inp_feat(416), I4 =>  inp_feat(269), I5 =>  inp_feat(341)); 
C_0_S_5_L_4_inst : LUT6 generic map(INIT => "1101011011011111110001111001111111011110100111011111111111111110") port map( O =>C_0_S_5_L_4_out, I0 =>  inp_feat(257), I1 =>  inp_feat(258), I2 =>  inp_feat(477), I3 =>  inp_feat(136), I4 =>  inp_feat(50), I5 =>  inp_feat(158)); 
C_0_S_5_L_5_inst : LUT6 generic map(INIT => "0010011010011101110101111101011110111011001111011111111111111001") port map( O =>C_0_S_5_L_5_out, I0 =>  inp_feat(257), I1 =>  inp_feat(334), I2 =>  inp_feat(477), I3 =>  inp_feat(136), I4 =>  inp_feat(50), I5 =>  inp_feat(158)); 
C_1_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111110111111001110000011101110111111001100100010000000") port map( O =>C_1_S_0_L_0_out, I0 =>  inp_feat(253), I1 =>  inp_feat(82), I2 =>  inp_feat(0), I3 =>  inp_feat(71), I4 =>  inp_feat(102), I5 =>  inp_feat(327)); 
C_1_S_0_L_1_inst : LUT6 generic map(INIT => "1111100110100010101011001110001111000001101100100000010010110001") port map( O =>C_1_S_0_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(445), I2 =>  inp_feat(29), I3 =>  inp_feat(58), I4 =>  inp_feat(373), I5 =>  inp_feat(431)); 
C_1_S_0_L_2_inst : LUT6 generic map(INIT => "1000111110001110000111010000000000000010101001000010100000000000") port map( O =>C_1_S_0_L_2_out, I0 =>  inp_feat(184), I1 =>  inp_feat(22), I2 =>  inp_feat(241), I3 =>  inp_feat(170), I4 =>  inp_feat(159), I5 =>  inp_feat(339)); 
C_1_S_0_L_3_inst : LUT6 generic map(INIT => "0100000010001010101000100000000011101110111000001110011010000000") port map( O =>C_1_S_0_L_3_out, I0 =>  inp_feat(71), I1 =>  inp_feat(74), I2 =>  inp_feat(72), I3 =>  inp_feat(315), I4 =>  inp_feat(325), I5 =>  inp_feat(354)); 
C_1_S_0_L_4_inst : LUT6 generic map(INIT => "1111101100001011100010100011010100110011000100110010001000101011") port map( O =>C_1_S_0_L_4_out, I0 =>  inp_feat(234), I1 =>  inp_feat(21), I2 =>  inp_feat(484), I3 =>  inp_feat(429), I4 =>  inp_feat(74), I5 =>  inp_feat(71)); 
C_1_S_0_L_5_inst : LUT6 generic map(INIT => "1111010101110101011100110111001100000000010001110101010111011111") port map( O =>C_1_S_0_L_5_out, I0 =>  inp_feat(458), I1 =>  inp_feat(387), I2 =>  inp_feat(237), I3 =>  inp_feat(481), I4 =>  inp_feat(73), I5 =>  inp_feat(177)); 
C_1_S_1_L_0_inst : LUT6 generic map(INIT => "1111100110100010101011001110001111000001101100100000010010110001") port map( O =>C_1_S_1_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(445), I2 =>  inp_feat(29), I3 =>  inp_feat(58), I4 =>  inp_feat(373), I5 =>  inp_feat(431)); 
C_1_S_1_L_1_inst : LUT6 generic map(INIT => "1000111110001110000111010000000000000010101001000010100000000000") port map( O =>C_1_S_1_L_1_out, I0 =>  inp_feat(184), I1 =>  inp_feat(22), I2 =>  inp_feat(241), I3 =>  inp_feat(170), I4 =>  inp_feat(159), I5 =>  inp_feat(339)); 
C_1_S_1_L_2_inst : LUT6 generic map(INIT => "0100000010001010101000100000000011101110111000001110011010000000") port map( O =>C_1_S_1_L_2_out, I0 =>  inp_feat(71), I1 =>  inp_feat(74), I2 =>  inp_feat(72), I3 =>  inp_feat(315), I4 =>  inp_feat(325), I5 =>  inp_feat(354)); 
C_1_S_1_L_3_inst : LUT6 generic map(INIT => "1111101100001011100010100011010100110011000100110010001000101011") port map( O =>C_1_S_1_L_3_out, I0 =>  inp_feat(234), I1 =>  inp_feat(21), I2 =>  inp_feat(484), I3 =>  inp_feat(429), I4 =>  inp_feat(74), I5 =>  inp_feat(71)); 
C_1_S_1_L_4_inst : LUT6 generic map(INIT => "1111010101110101011100110111001100000000010001110101010111011111") port map( O =>C_1_S_1_L_4_out, I0 =>  inp_feat(458), I1 =>  inp_feat(387), I2 =>  inp_feat(237), I3 =>  inp_feat(481), I4 =>  inp_feat(73), I5 =>  inp_feat(177)); 
C_1_S_1_L_5_inst : LUT6 generic map(INIT => "0000100001001101101011000000110100100011111111100000101000000010") port map( O =>C_1_S_1_L_5_out, I0 =>  inp_feat(413), I1 =>  inp_feat(315), I2 =>  inp_feat(127), I3 =>  inp_feat(410), I4 =>  inp_feat(29), I5 =>  inp_feat(161)); 
C_1_S_2_L_0_inst : LUT6 generic map(INIT => "1011101010111011111111111111111010111110111000001111111011010000") port map( O =>C_1_S_2_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(157), I2 =>  inp_feat(277), I3 =>  inp_feat(321), I4 =>  inp_feat(395), I5 =>  inp_feat(241)); 
C_1_S_2_L_1_inst : LUT6 generic map(INIT => "0001010000100000001100101010001010111100000000001111111010100000") port map( O =>C_1_S_2_L_1_out, I0 =>  inp_feat(170), I1 =>  inp_feat(379), I2 =>  inp_feat(234), I3 =>  inp_feat(0), I4 =>  inp_feat(356), I5 =>  inp_feat(287)); 
C_1_S_2_L_2_inst : LUT6 generic map(INIT => "1110111010111000111010000010100001110010110000000000000000000000") port map( O =>C_1_S_2_L_2_out, I0 =>  inp_feat(180), I1 =>  inp_feat(58), I2 =>  inp_feat(234), I3 =>  inp_feat(319), I4 =>  inp_feat(74), I5 =>  inp_feat(315)); 
C_1_S_2_L_3_inst : LUT6 generic map(INIT => "0111101001100100100010001100000000001110110011001110000000000000") port map( O =>C_1_S_2_L_3_out, I0 =>  inp_feat(180), I1 =>  inp_feat(15), I2 =>  inp_feat(319), I3 =>  inp_feat(170), I4 =>  inp_feat(410), I5 =>  inp_feat(164)); 
C_1_S_2_L_4_inst : LUT6 generic map(INIT => "1011110110000001101011001101000011010101010101011100000000000000") port map( O =>C_1_S_2_L_4_out, I0 =>  inp_feat(182), I1 =>  inp_feat(410), I2 =>  inp_feat(82), I3 =>  inp_feat(52), I4 =>  inp_feat(346), I5 =>  inp_feat(379)); 
C_1_S_2_L_5_inst : LUT6 generic map(INIT => "0000101000100000110000110010000011101110110010001101111110000000") port map( O =>C_1_S_2_L_5_out, I0 =>  inp_feat(164), I1 =>  inp_feat(52), I2 =>  inp_feat(277), I3 =>  inp_feat(177), I4 =>  inp_feat(173), I5 =>  inp_feat(38)); 
C_1_S_3_L_0_inst : LUT6 generic map(INIT => "0010101010110010110000110010001101011010110100001000001000000000") port map( O =>C_1_S_3_L_0_out, I0 =>  inp_feat(347), I1 =>  inp_feat(24), I2 =>  inp_feat(159), I3 =>  inp_feat(170), I4 =>  inp_feat(410), I5 =>  inp_feat(164)); 
C_1_S_3_L_1_inst : LUT6 generic map(INIT => "1001000110010011110110111001001010111111101100111101000000010000") port map( O =>C_1_S_3_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(373), I2 =>  inp_feat(15), I3 =>  inp_feat(159), I4 =>  inp_feat(325), I5 =>  inp_feat(354)); 
C_1_S_3_L_2_inst : LUT6 generic map(INIT => "1010010111100111110011001110101010000100111111000000100010101000") port map( O =>C_1_S_3_L_2_out, I0 =>  inp_feat(296), I1 =>  inp_feat(74), I2 =>  inp_feat(103), I3 =>  inp_feat(395), I4 =>  inp_feat(29), I5 =>  inp_feat(410)); 
C_1_S_3_L_3_inst : LUT6 generic map(INIT => "1110111001001110110011100111111100001011000111111100111011111111") port map( O =>C_1_S_3_L_3_out, I0 =>  inp_feat(336), I1 =>  inp_feat(454), I2 =>  inp_feat(17), I3 =>  inp_feat(291), I4 =>  inp_feat(221), I5 =>  inp_feat(96)); 
C_1_S_3_L_4_inst : LUT6 generic map(INIT => "0010111100010101110111110100000011111111010011010111001001110100") port map( O =>C_1_S_3_L_4_out, I0 =>  inp_feat(227), I1 =>  inp_feat(283), I2 =>  inp_feat(479), I3 =>  inp_feat(180), I4 =>  inp_feat(419), I5 =>  inp_feat(179)); 
C_1_S_3_L_5_inst : LUT6 generic map(INIT => "1100111011001000100010001111101001111011111110000000101010001010") port map( O =>C_1_S_3_L_5_out, I0 =>  inp_feat(234), I1 =>  inp_feat(71), I2 =>  inp_feat(474), I3 =>  inp_feat(221), I4 =>  inp_feat(361), I5 =>  inp_feat(126)); 
C_1_S_4_L_0_inst : LUT6 generic map(INIT => "1110001100001100001000100100111001101100000011000001001011111111") port map( O =>C_1_S_4_L_0_out, I0 =>  inp_feat(205), I1 =>  inp_feat(10), I2 =>  inp_feat(194), I3 =>  inp_feat(420), I4 =>  inp_feat(170), I5 =>  inp_feat(490)); 
C_1_S_4_L_1_inst : LUT6 generic map(INIT => "0001011100101000001111101111010010111111111111111111101010110100") port map( O =>C_1_S_4_L_1_out, I0 =>  inp_feat(508), I1 =>  inp_feat(445), I2 =>  inp_feat(241), I3 =>  inp_feat(7), I4 =>  inp_feat(461), I5 =>  inp_feat(282)); 
C_1_S_4_L_2_inst : LUT6 generic map(INIT => "1110100011001100011011101110110000011111000100111110111100111101") port map( O =>C_1_S_4_L_2_out, I0 =>  inp_feat(476), I1 =>  inp_feat(122), I2 =>  inp_feat(181), I3 =>  inp_feat(0), I4 =>  inp_feat(330), I5 =>  inp_feat(398)); 
C_1_S_4_L_3_inst : LUT6 generic map(INIT => "0011111011111111001111011111101100101001111110000100000011000000") port map( O =>C_1_S_4_L_3_out, I0 =>  inp_feat(483), I1 =>  inp_feat(392), I2 =>  inp_feat(277), I3 =>  inp_feat(395), I4 =>  inp_feat(410), I5 =>  inp_feat(164)); 
C_1_S_4_L_4_inst : LUT6 generic map(INIT => "0111111011001110010110011111111111101111111111010000111111111111") port map( O =>C_1_S_4_L_4_out, I0 =>  inp_feat(21), I1 =>  inp_feat(419), I2 =>  inp_feat(196), I3 =>  inp_feat(356), I4 =>  inp_feat(60), I5 =>  inp_feat(181)); 
C_1_S_4_L_5_inst : LUT6 generic map(INIT => "1111110111111001110100010000000111111111111101111111101100011011") port map( O =>C_1_S_4_L_5_out, I0 =>  inp_feat(127), I1 =>  inp_feat(348), I2 =>  inp_feat(71), I3 =>  inp_feat(173), I4 =>  inp_feat(120), I5 =>  inp_feat(38)); 
C_1_S_5_L_0_inst : LUT6 generic map(INIT => "1000100010010100000011101111100000110010110100100000100111001111") port map( O =>C_1_S_5_L_0_out, I0 =>  inp_feat(484), I1 =>  inp_feat(56), I2 =>  inp_feat(343), I3 =>  inp_feat(420), I4 =>  inp_feat(170), I5 =>  inp_feat(490)); 
C_1_S_5_L_1_inst : LUT6 generic map(INIT => "0111110010101110000000001010001000110110111111001000000011000000") port map( O =>C_1_S_5_L_1_out, I0 =>  inp_feat(71), I1 =>  inp_feat(153), I2 =>  inp_feat(319), I3 =>  inp_feat(318), I4 =>  inp_feat(74), I5 =>  inp_feat(242)); 
C_1_S_5_L_2_inst : LUT6 generic map(INIT => "0010001000100000001100110001111111111111110101111110111101101011") port map( O =>C_1_S_5_L_2_out, I0 =>  inp_feat(205), I1 =>  inp_feat(179), I2 =>  inp_feat(59), I3 =>  inp_feat(60), I4 =>  inp_feat(307), I5 =>  inp_feat(46)); 
C_1_S_5_L_3_inst : LUT6 generic map(INIT => "1101110011001000011011010001000111101111111110010011100111111111") port map( O =>C_1_S_5_L_3_out, I0 =>  inp_feat(428), I1 =>  inp_feat(96), I2 =>  inp_feat(384), I3 =>  inp_feat(175), I4 =>  inp_feat(205), I5 =>  inp_feat(38)); 
C_1_S_5_L_4_inst : LUT6 generic map(INIT => "0000001010110011010011001110110011101100111111110000000011111010") port map( O =>C_1_S_5_L_4_out, I0 =>  inp_feat(178), I1 =>  inp_feat(231), I2 =>  inp_feat(93), I3 =>  inp_feat(77), I4 =>  inp_feat(244), I5 =>  inp_feat(412)); 
C_1_S_5_L_5_inst : LUT6 generic map(INIT => "1101110111111111111111111110111000111110110011101100101110001100") port map( O =>C_1_S_5_L_5_out, I0 =>  inp_feat(158), I1 =>  inp_feat(385), I2 =>  inp_feat(443), I3 =>  inp_feat(50), I4 =>  inp_feat(504), I5 =>  inp_feat(87)); 
C_2_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111111110100011111101111010001110110010000000") port map( O =>C_2_S_0_L_0_out, I0 =>  inp_feat(315), I1 =>  inp_feat(432), I2 =>  inp_feat(435), I3 =>  inp_feat(0), I4 =>  inp_feat(102), I5 =>  inp_feat(58)); 
C_2_S_0_L_1_inst : LUT6 generic map(INIT => "1111101111010001000001100001011000010010001011100001111100001100") port map( O =>C_2_S_0_L_1_out, I0 =>  inp_feat(371), I1 =>  inp_feat(244), I2 =>  inp_feat(204), I3 =>  inp_feat(159), I4 =>  inp_feat(71), I5 =>  inp_feat(180)); 
C_2_S_0_L_2_inst : LUT6 generic map(INIT => "1110101110101010101111110110110000011100101111011110110011001100") port map( O =>C_2_S_0_L_2_out, I0 =>  inp_feat(292), I1 =>  inp_feat(351), I2 =>  inp_feat(313), I3 =>  inp_feat(279), I4 =>  inp_feat(378), I5 =>  inp_feat(159)); 
C_2_S_0_L_3_inst : LUT6 generic map(INIT => "0001000010011000100110001000000011111111111011001111110011010000") port map( O =>C_2_S_0_L_3_out, I0 =>  inp_feat(189), I1 =>  inp_feat(71), I2 =>  inp_feat(82), I3 =>  inp_feat(159), I4 =>  inp_feat(180), I5 =>  inp_feat(421)); 
C_2_S_0_L_4_inst : LUT6 generic map(INIT => "1111111101110111111111011111101101110100011101001111111111111100") port map( O =>C_2_S_0_L_4_out, I0 =>  inp_feat(126), I1 =>  inp_feat(80), I2 =>  inp_feat(227), I3 =>  inp_feat(505), I4 =>  inp_feat(39), I5 =>  inp_feat(190)); 
C_2_S_0_L_5_inst : LUT6 generic map(INIT => "1010001110001111000100011100111111101111111100101111111101101111") port map( O =>C_2_S_0_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(242), I2 =>  inp_feat(194), I3 =>  inp_feat(75), I4 =>  inp_feat(227), I5 =>  inp_feat(39)); 
C_2_S_1_L_0_inst : LUT6 generic map(INIT => "1111101111010001000001100001011000010010001011100001111100001100") port map( O =>C_2_S_1_L_0_out, I0 =>  inp_feat(371), I1 =>  inp_feat(244), I2 =>  inp_feat(204), I3 =>  inp_feat(159), I4 =>  inp_feat(71), I5 =>  inp_feat(180)); 
C_2_S_1_L_1_inst : LUT6 generic map(INIT => "1110101110101010101111110110110000011100101111011110110011001100") port map( O =>C_2_S_1_L_1_out, I0 =>  inp_feat(292), I1 =>  inp_feat(351), I2 =>  inp_feat(313), I3 =>  inp_feat(279), I4 =>  inp_feat(378), I5 =>  inp_feat(159)); 
C_2_S_1_L_2_inst : LUT6 generic map(INIT => "0001000010011000100110001000000011111111111011001111110011010000") port map( O =>C_2_S_1_L_2_out, I0 =>  inp_feat(189), I1 =>  inp_feat(71), I2 =>  inp_feat(82), I3 =>  inp_feat(159), I4 =>  inp_feat(180), I5 =>  inp_feat(421)); 
C_2_S_1_L_3_inst : LUT6 generic map(INIT => "1111111101110111111111011111101101110100011101001111111111111100") port map( O =>C_2_S_1_L_3_out, I0 =>  inp_feat(126), I1 =>  inp_feat(80), I2 =>  inp_feat(227), I3 =>  inp_feat(505), I4 =>  inp_feat(39), I5 =>  inp_feat(190)); 
C_2_S_1_L_4_inst : LUT6 generic map(INIT => "1010001110001111000100011100111111101111111100101111111101101111") port map( O =>C_2_S_1_L_4_out, I0 =>  inp_feat(82), I1 =>  inp_feat(242), I2 =>  inp_feat(194), I3 =>  inp_feat(75), I4 =>  inp_feat(227), I5 =>  inp_feat(39)); 
C_2_S_1_L_5_inst : LUT6 generic map(INIT => "1010000010101100111000111010100000000100111001001111111110000000") port map( O =>C_2_S_1_L_5_out, I0 =>  inp_feat(159), I1 =>  inp_feat(253), I2 =>  inp_feat(296), I3 =>  inp_feat(287), I4 =>  inp_feat(320), I5 =>  inp_feat(26)); 
C_2_S_2_L_0_inst : LUT6 generic map(INIT => "1000100110001111100000111110101011101111101111111110111101000010") port map( O =>C_2_S_2_L_0_out, I0 =>  inp_feat(472), I1 =>  inp_feat(74), I2 =>  inp_feat(312), I3 =>  inp_feat(326), I4 =>  inp_feat(420), I5 =>  inp_feat(363)); 
C_2_S_2_L_1_inst : LUT6 generic map(INIT => "0111110111110011001010111111111100110111001011100001111100011101") port map( O =>C_2_S_2_L_1_out, I0 =>  inp_feat(91), I1 =>  inp_feat(306), I2 =>  inp_feat(111), I3 =>  inp_feat(120), I4 =>  inp_feat(315), I5 =>  inp_feat(325)); 
C_2_S_2_L_2_inst : LUT6 generic map(INIT => "1011110110010001001111011011111111111111111011001011111110100010") port map( O =>C_2_S_2_L_2_out, I0 =>  inp_feat(489), I1 =>  inp_feat(368), I2 =>  inp_feat(481), I3 =>  inp_feat(454), I4 =>  inp_feat(22), I5 =>  inp_feat(363)); 
C_2_S_2_L_3_inst : LUT6 generic map(INIT => "0010101111010000001011101111101111101110111010101100111010100010") port map( O =>C_2_S_2_L_3_out, I0 =>  inp_feat(315), I1 =>  inp_feat(128), I2 =>  inp_feat(210), I3 =>  inp_feat(420), I4 =>  inp_feat(341), I5 =>  inp_feat(363)); 
C_2_S_2_L_4_inst : LUT6 generic map(INIT => "1101101110100010101111111111111000010011001000111110110101001100") port map( O =>C_2_S_2_L_4_out, I0 =>  inp_feat(209), I1 =>  inp_feat(289), I2 =>  inp_feat(451), I3 =>  inp_feat(243), I4 =>  inp_feat(458), I5 =>  inp_feat(315)); 
C_2_S_2_L_5_inst : LUT6 generic map(INIT => "0001110011011010000110111000111111111111111111111010110111111111") port map( O =>C_2_S_2_L_5_out, I0 =>  inp_feat(305), I1 =>  inp_feat(379), I2 =>  inp_feat(225), I3 =>  inp_feat(257), I4 =>  inp_feat(164), I5 =>  inp_feat(372)); 
C_2_S_3_L_0_inst : LUT6 generic map(INIT => "0111110000110101100011000110110011111111111111011110011011111111") port map( O =>C_2_S_3_L_0_out, I0 =>  inp_feat(282), I1 =>  inp_feat(423), I2 =>  inp_feat(38), I3 =>  inp_feat(253), I4 =>  inp_feat(391), I5 =>  inp_feat(320)); 
C_2_S_3_L_1_inst : LUT6 generic map(INIT => "1010100001001110110000001110100011111111111111111111111110000000") port map( O =>C_2_S_3_L_1_out, I0 =>  inp_feat(159), I1 =>  inp_feat(234), I2 =>  inp_feat(267), I3 =>  inp_feat(196), I4 =>  inp_feat(243), I5 =>  inp_feat(246)); 
C_2_S_3_L_2_inst : LUT6 generic map(INIT => "1010000011000100111111011010011000101000111010000110111011000000") port map( O =>C_2_S_3_L_2_out, I0 =>  inp_feat(315), I1 =>  inp_feat(153), I2 =>  inp_feat(319), I3 =>  inp_feat(405), I4 =>  inp_feat(84), I5 =>  inp_feat(190)); 
C_2_S_3_L_3_inst : LUT6 generic map(INIT => "1000111111100111001101101110111101001111111111100110101011111100") port map( O =>C_2_S_3_L_3_out, I0 =>  inp_feat(432), I1 =>  inp_feat(136), I2 =>  inp_feat(343), I3 =>  inp_feat(289), I4 =>  inp_feat(151), I5 =>  inp_feat(399)); 
C_2_S_3_L_4_inst : LUT6 generic map(INIT => "1011111010111110000011001110001011111110111010101111101010100000") port map( O =>C_2_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(234), I2 =>  inp_feat(459), I3 =>  inp_feat(461), I4 =>  inp_feat(82), I5 =>  inp_feat(158)); 
C_2_S_3_L_5_inst : LUT6 generic map(INIT => "0111111110111111111111111111001001110011101110101011000011110000") port map( O =>C_2_S_3_L_5_out, I0 =>  inp_feat(488), I1 =>  inp_feat(301), I2 =>  inp_feat(444), I3 =>  inp_feat(296), I4 =>  inp_feat(99), I5 =>  inp_feat(201)); 
C_2_S_4_L_0_inst : LUT6 generic map(INIT => "1100100000101010111010101110101111101000001011110011011100011111") port map( O =>C_2_S_4_L_0_out, I0 =>  inp_feat(74), I1 =>  inp_feat(164), I2 =>  inp_feat(174), I3 =>  inp_feat(13), I4 =>  inp_feat(218), I5 =>  inp_feat(505)); 
C_2_S_4_L_1_inst : LUT6 generic map(INIT => "1011110100111110000111100011111111111111111111101111110100101110") port map( O =>C_2_S_4_L_1_out, I0 =>  inp_feat(56), I1 =>  inp_feat(378), I2 =>  inp_feat(232), I3 =>  inp_feat(153), I4 =>  inp_feat(420), I5 =>  inp_feat(289)); 
C_2_S_4_L_2_inst : LUT6 generic map(INIT => "1101101111101111111001011111110000000000111111101111110101101001") port map( O =>C_2_S_4_L_2_out, I0 =>  inp_feat(415), I1 =>  inp_feat(335), I2 =>  inp_feat(68), I3 =>  inp_feat(240), I4 =>  inp_feat(83), I5 =>  inp_feat(108)); 
C_2_S_4_L_3_inst : LUT6 generic map(INIT => "1111100110011111111010001111111100110011000010111111111100001000") port map( O =>C_2_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(257), I2 =>  inp_feat(338), I3 =>  inp_feat(74), I4 =>  inp_feat(481), I5 =>  inp_feat(82)); 
C_2_S_4_L_4_inst : LUT6 generic map(INIT => "0011110100101101101001111001101011101010101010000010100000001010") port map( O =>C_2_S_4_L_4_out, I0 =>  inp_feat(234), I1 =>  inp_feat(341), I2 =>  inp_feat(363), I3 =>  inp_feat(460), I4 =>  inp_feat(205), I5 =>  inp_feat(134)); 
C_2_S_4_L_5_inst : LUT6 generic map(INIT => "1101111010000000110010100111100011101110101000100110110001100000") port map( O =>C_2_S_4_L_5_out, I0 =>  inp_feat(71), I1 =>  inp_feat(379), I2 =>  inp_feat(82), I3 =>  inp_feat(292), I4 =>  inp_feat(205), I5 =>  inp_feat(134)); 
C_2_S_5_L_0_inst : LUT6 generic map(INIT => "1010111111111111111111101111111110001000111111001111111100111111") port map( O =>C_2_S_5_L_0_out, I0 =>  inp_feat(399), I1 =>  inp_feat(344), I2 =>  inp_feat(373), I3 =>  inp_feat(380), I4 =>  inp_feat(83), I5 =>  inp_feat(182)); 
C_2_S_5_L_1_inst : LUT6 generic map(INIT => "0000001001011110111001100101111100101000010011111101110011111111") port map( O =>C_2_S_5_L_1_out, I0 =>  inp_feat(71), I1 =>  inp_feat(164), I2 =>  inp_feat(460), I3 =>  inp_feat(489), I4 =>  inp_feat(257), I5 =>  inp_feat(267)); 
C_2_S_5_L_2_inst : LUT6 generic map(INIT => "1011000011011110111011001110110000101110111110110010100001101110") port map( O =>C_2_S_5_L_2_out, I0 =>  inp_feat(71), I1 =>  inp_feat(234), I2 =>  inp_feat(6), I3 =>  inp_feat(257), I4 =>  inp_feat(243), I5 =>  inp_feat(267)); 
C_2_S_5_L_3_inst : LUT6 generic map(INIT => "0001110100011101010111010011111111101111111011110110111011111110") port map( O =>C_2_S_5_L_3_out, I0 =>  inp_feat(133), I1 =>  inp_feat(467), I2 =>  inp_feat(306), I3 =>  inp_feat(280), I4 =>  inp_feat(82), I5 =>  inp_feat(92)); 
C_2_S_5_L_4_inst : LUT6 generic map(INIT => "0101111011111110100010101110010011111110111011001111110011000000") port map( O =>C_2_S_5_L_4_out, I0 =>  inp_feat(234), I1 =>  inp_feat(0), I2 =>  inp_feat(459), I3 =>  inp_feat(461), I4 =>  inp_feat(82), I5 =>  inp_feat(158)); 
C_2_S_5_L_5_inst : LUT6 generic map(INIT => "1110011111110111100110111011111100001101011111110010100111101111") port map( O =>C_2_S_5_L_5_out, I0 =>  inp_feat(478), I1 =>  inp_feat(234), I2 =>  inp_feat(440), I3 =>  inp_feat(320), I4 =>  inp_feat(31), I5 =>  inp_feat(296)); 
C_3_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111101010000011101100111010001110000010000000") port map( O =>C_3_S_0_L_0_out, I0 =>  inp_feat(71), I1 =>  inp_feat(436), I2 =>  inp_feat(82), I3 =>  inp_feat(0), I4 =>  inp_feat(102), I5 =>  inp_feat(327)); 
C_3_S_0_L_1_inst : LUT6 generic map(INIT => "1111101110110010111100100001001000010111101000111101100111111011") port map( O =>C_3_S_0_L_1_out, I0 =>  inp_feat(319), I1 =>  inp_feat(257), I2 =>  inp_feat(15), I3 =>  inp_feat(159), I4 =>  inp_feat(325), I5 =>  inp_feat(497)); 
C_3_S_0_L_2_inst : LUT6 generic map(INIT => "1001010100010001010011010101111111111011111111011110111011110111") port map( O =>C_3_S_0_L_2_out, I0 =>  inp_feat(116), I1 =>  inp_feat(153), I2 =>  inp_feat(394), I3 =>  inp_feat(194), I4 =>  inp_feat(346), I5 =>  inp_feat(84)); 
C_3_S_0_L_3_inst : LUT6 generic map(INIT => "0111111011011000110011000000000011110110111100011110100010000000") port map( O =>C_3_S_0_L_3_out, I0 =>  inp_feat(29), I1 =>  inp_feat(74), I2 =>  inp_feat(253), I3 =>  inp_feat(159), I4 =>  inp_feat(0), I5 =>  inp_feat(434)); 
C_3_S_0_L_4_inst : LUT6 generic map(INIT => "0000110010001111010011001111111111101010110010101110100011101100") port map( O =>C_3_S_0_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(325), I2 =>  inp_feat(102), I3 =>  inp_feat(257), I4 =>  inp_feat(404), I5 =>  inp_feat(386)); 
C_3_S_0_L_5_inst : LUT6 generic map(INIT => "1101111110111111110110101111111001100111011011001011011011101011") port map( O =>C_3_S_0_L_5_out, I0 =>  inp_feat(474), I1 =>  inp_feat(319), I2 =>  inp_feat(370), I3 =>  inp_feat(83), I4 =>  inp_feat(95), I5 =>  inp_feat(407)); 
C_3_S_1_L_0_inst : LUT6 generic map(INIT => "1111101110110010111100100001001000010111101000111101100111111011") port map( O =>C_3_S_1_L_0_out, I0 =>  inp_feat(319), I1 =>  inp_feat(257), I2 =>  inp_feat(15), I3 =>  inp_feat(159), I4 =>  inp_feat(325), I5 =>  inp_feat(497)); 
C_3_S_1_L_1_inst : LUT6 generic map(INIT => "1001010100010001010011010101111111111011111111011110111011110111") port map( O =>C_3_S_1_L_1_out, I0 =>  inp_feat(116), I1 =>  inp_feat(153), I2 =>  inp_feat(394), I3 =>  inp_feat(194), I4 =>  inp_feat(346), I5 =>  inp_feat(84)); 
C_3_S_1_L_2_inst : LUT6 generic map(INIT => "0111111011011000110011000000000011110110111100011110100010000000") port map( O =>C_3_S_1_L_2_out, I0 =>  inp_feat(29), I1 =>  inp_feat(74), I2 =>  inp_feat(253), I3 =>  inp_feat(159), I4 =>  inp_feat(0), I5 =>  inp_feat(434)); 
C_3_S_1_L_3_inst : LUT6 generic map(INIT => "0000110010001111010011001111111111101010110010101110100011101100") port map( O =>C_3_S_1_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(325), I2 =>  inp_feat(102), I3 =>  inp_feat(257), I4 =>  inp_feat(404), I5 =>  inp_feat(386)); 
C_3_S_1_L_4_inst : LUT6 generic map(INIT => "1101111110111111110110101111111001100111011011001011011011101011") port map( O =>C_3_S_1_L_4_out, I0 =>  inp_feat(474), I1 =>  inp_feat(319), I2 =>  inp_feat(370), I3 =>  inp_feat(83), I4 =>  inp_feat(95), I5 =>  inp_feat(407)); 
C_3_S_1_L_5_inst : LUT6 generic map(INIT => "1111001110110011000100111111111100000001010100100101000111110111") port map( O =>C_3_S_1_L_5_out, I0 =>  inp_feat(59), I1 =>  inp_feat(111), I2 =>  inp_feat(323), I3 =>  inp_feat(1), I4 =>  inp_feat(251), I5 =>  inp_feat(29)); 
C_3_S_2_L_0_inst : LUT6 generic map(INIT => "0110011011100000010111000000000011111111010011101011111111001110") port map( O =>C_3_S_2_L_0_out, I0 =>  inp_feat(180), I1 =>  inp_feat(170), I2 =>  inp_feat(451), I3 =>  inp_feat(159), I4 =>  inp_feat(346), I5 =>  inp_feat(84)); 
C_3_S_2_L_1_inst : LUT6 generic map(INIT => "1110111011011000101011001000000011111110111110001110000010000000") port map( O =>C_3_S_2_L_1_out, I0 =>  inp_feat(455), I1 =>  inp_feat(74), I2 =>  inp_feat(190), I3 =>  inp_feat(159), I4 =>  inp_feat(0), I5 =>  inp_feat(434)); 
C_3_S_2_L_2_inst : LUT6 generic map(INIT => "0100011010011000011010001100000011111010111010001010100000100000") port map( O =>C_3_S_2_L_2_out, I0 =>  inp_feat(71), I1 =>  inp_feat(464), I2 =>  inp_feat(234), I3 =>  inp_feat(74), I4 =>  inp_feat(228), I5 =>  inp_feat(434)); 
C_3_S_2_L_3_inst : LUT6 generic map(INIT => "1101010001011100111111111111110111110111111111111111111111110110") port map( O =>C_3_S_2_L_3_out, I0 =>  inp_feat(372), I1 =>  inp_feat(210), I2 =>  inp_feat(160), I3 =>  inp_feat(326), I4 =>  inp_feat(195), I5 =>  inp_feat(386)); 
C_3_S_2_L_4_inst : LUT6 generic map(INIT => "0111111101101110111111110101110111101111111111110011111101011111") port map( O =>C_3_S_2_L_4_out, I0 =>  inp_feat(195), I1 =>  inp_feat(73), I2 =>  inp_feat(361), I3 =>  inp_feat(492), I4 =>  inp_feat(420), I5 =>  inp_feat(202)); 
C_3_S_2_L_5_inst : LUT6 generic map(INIT => "1110111011111101111001000111111100001100111111110000100000001110") port map( O =>C_3_S_2_L_5_out, I0 =>  inp_feat(230), I1 =>  inp_feat(253), I2 =>  inp_feat(45), I3 =>  inp_feat(419), I4 =>  inp_feat(29), I5 =>  inp_feat(410)); 
C_3_S_3_L_0_inst : LUT6 generic map(INIT => "0101110101011100010111010100000011011111110111001101000100010000") port map( O =>C_3_S_3_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(253), I2 =>  inp_feat(190), I3 =>  inp_feat(159), I4 =>  inp_feat(0), I5 =>  inp_feat(434)); 
C_3_S_3_L_1_inst : LUT6 generic map(INIT => "1001000101000001111110110111111100010101111011110011111011110010") port map( O =>C_3_S_3_L_1_out, I0 =>  inp_feat(215), I1 =>  inp_feat(0), I2 =>  inp_feat(288), I3 =>  inp_feat(378), I4 =>  inp_feat(168), I5 =>  inp_feat(72)); 
C_3_S_3_L_2_inst : LUT6 generic map(INIT => "1111101110111011101101110111101101000011011000101110111010000000") port map( O =>C_3_S_3_L_2_out, I0 =>  inp_feat(74), I1 =>  inp_feat(279), I2 =>  inp_feat(234), I3 =>  inp_feat(0), I4 =>  inp_feat(356), I5 =>  inp_feat(72)); 
C_3_S_3_L_3_inst : LUT6 generic map(INIT => "0101011110000100111010101110000011111111101011001111111001101010") port map( O =>C_3_S_3_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(234), I2 =>  inp_feat(464), I3 =>  inp_feat(74), I4 =>  inp_feat(228), I5 =>  inp_feat(434)); 
C_3_S_3_L_4_inst : LUT6 generic map(INIT => "1010110011101111001111100111111100101000110111111111110111111110") port map( O =>C_3_S_3_L_4_out, I0 =>  inp_feat(29), I1 =>  inp_feat(315), I2 =>  inp_feat(102), I3 =>  inp_feat(91), I4 =>  inp_feat(122), I5 =>  inp_feat(242)); 
C_3_S_3_L_5_inst : LUT6 generic map(INIT => "0001110101000110000111000011000111100110001000101111111111111011") port map( O =>C_3_S_3_L_5_out, I0 =>  inp_feat(307), I1 =>  inp_feat(486), I2 =>  inp_feat(505), I3 =>  inp_feat(190), I4 =>  inp_feat(199), I5 =>  inp_feat(111)); 
C_3_S_4_L_0_inst : LUT6 generic map(INIT => "0110110011000100101010010001111011101100111010001110111011000000") port map( O =>C_3_S_4_L_0_out, I0 =>  inp_feat(432), I1 =>  inp_feat(315), I2 =>  inp_feat(379), I3 =>  inp_feat(112), I4 =>  inp_feat(68), I5 =>  inp_feat(217)); 
C_3_S_4_L_1_inst : LUT6 generic map(INIT => "1101110010101000111011001010110000111000111100001111110000111100") port map( O =>C_3_S_4_L_1_out, I0 =>  inp_feat(253), I1 =>  inp_feat(52), I2 =>  inp_feat(346), I3 =>  inp_feat(191), I4 =>  inp_feat(128), I5 =>  inp_feat(21)); 
C_3_S_4_L_2_inst : LUT6 generic map(INIT => "0010010000010110000110101100111111100011111101111111111111111111") port map( O =>C_3_S_4_L_2_out, I0 =>  inp_feat(224), I1 =>  inp_feat(305), I2 =>  inp_feat(272), I3 =>  inp_feat(361), I4 =>  inp_feat(300), I5 =>  inp_feat(202)); 
C_3_S_4_L_3_inst : LUT6 generic map(INIT => "0100101000101111011011101110111111111110111111111000110011111111") port map( O =>C_3_S_4_L_3_out, I0 =>  inp_feat(395), I1 =>  inp_feat(373), I2 =>  inp_feat(226), I3 =>  inp_feat(242), I4 =>  inp_feat(306), I5 =>  inp_feat(355)); 
C_3_S_4_L_4_inst : LUT6 generic map(INIT => "1011001111101010010111110011111111111111111111110011001111111111") port map( O =>C_3_S_4_L_4_out, I0 =>  inp_feat(235), I1 =>  inp_feat(419), I2 =>  inp_feat(437), I3 =>  inp_feat(242), I4 =>  inp_feat(410), I5 =>  inp_feat(57)); 
C_3_S_4_L_5_inst : LUT6 generic map(INIT => "0001010100010111101010111111111011111111001111111001101111111011") port map( O =>C_3_S_4_L_5_out, I0 =>  inp_feat(488), I1 =>  inp_feat(419), I2 =>  inp_feat(393), I3 =>  inp_feat(220), I4 =>  inp_feat(269), I5 =>  inp_feat(57)); 
C_3_S_5_L_0_inst : LUT6 generic map(INIT => "0010001000101100101010001100000011101110111010001010100000001000") port map( O =>C_3_S_5_L_0_out, I0 =>  inp_feat(71), I1 =>  inp_feat(234), I2 =>  inp_feat(464), I3 =>  inp_feat(74), I4 =>  inp_feat(228), I5 =>  inp_feat(434)); 
C_3_S_5_L_1_inst : LUT6 generic map(INIT => "1111111101111110110101001101111111101100001011101101000011111101") port map( O =>C_3_S_5_L_1_out, I0 =>  inp_feat(1), I1 =>  inp_feat(61), I2 =>  inp_feat(489), I3 =>  inp_feat(251), I4 =>  inp_feat(277), I5 =>  inp_feat(118)); 
C_3_S_5_L_2_inst : LUT6 generic map(INIT => "0100010000001100011111000101111110101100111111111111101111110111") port map( O =>C_3_S_5_L_2_out, I0 =>  inp_feat(476), I1 =>  inp_feat(227), I2 =>  inp_feat(282), I3 =>  inp_feat(59), I4 =>  inp_feat(120), I5 =>  inp_feat(122)); 
C_3_S_5_L_3_inst : LUT6 generic map(INIT => "1111010100101111011010101111100111111111111111111111110111111111") port map( O =>C_3_S_5_L_3_out, I0 =>  inp_feat(96), I1 =>  inp_feat(13), I2 =>  inp_feat(407), I3 =>  inp_feat(128), I4 =>  inp_feat(68), I5 =>  inp_feat(217)); 
C_3_S_5_L_4_inst : LUT6 generic map(INIT => "1110110011111110011001101100111001101010000000100000000000101010") port map( O =>C_3_S_5_L_4_out, I0 =>  inp_feat(74), I1 =>  inp_feat(319), I2 =>  inp_feat(456), I3 =>  inp_feat(339), I4 =>  inp_feat(176), I5 =>  inp_feat(190)); 
C_3_S_5_L_5_inst : LUT6 generic map(INIT => "0010100110101010011001100110001111111111111101011111111110000001") port map( O =>C_3_S_5_L_5_out, I0 =>  inp_feat(403), I1 =>  inp_feat(277), I2 =>  inp_feat(226), I3 =>  inp_feat(44), I4 =>  inp_feat(39), I5 =>  inp_feat(355)); 
C_4_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111011101100000011111110111010001110000000000000") port map( O =>C_4_S_0_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(58), I2 =>  inp_feat(82), I3 =>  inp_feat(0), I4 =>  inp_feat(102), I5 =>  inp_feat(327)); 
C_4_S_0_L_1_inst : LUT6 generic map(INIT => "0000010111001110110011101100000011111111111011111100111011000000") port map( O =>C_4_S_0_L_1_out, I0 =>  inp_feat(405), I1 =>  inp_feat(494), I2 =>  inp_feat(444), I3 =>  inp_feat(28), I4 =>  inp_feat(222), I5 =>  inp_feat(312)); 
C_4_S_0_L_2_inst : LUT6 generic map(INIT => "1111111001111100111111000110000011111100011011001110000010000000") port map( O =>C_4_S_0_L_2_out, I0 =>  inp_feat(153), I1 =>  inp_feat(435), I2 =>  inp_feat(71), I3 =>  inp_feat(55), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_0_L_3_inst : LUT6 generic map(INIT => "0111010111111110111111001010100001111111011010001110100000000000") port map( O =>C_4_S_0_L_3_out, I0 =>  inp_feat(234), I1 =>  inp_feat(464), I2 =>  inp_feat(315), I3 =>  inp_feat(71), I4 =>  inp_feat(74), I5 =>  inp_feat(82)); 
C_4_S_0_L_4_inst : LUT6 generic map(INIT => "1111111111101010111111100110100011101010110010001111100010000000") port map( O =>C_4_S_0_L_4_out, I0 =>  inp_feat(159), I1 =>  inp_feat(432), I2 =>  inp_feat(71), I3 =>  inp_feat(0), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_0_L_5_inst : LUT6 generic map(INIT => "1101110111111110011110101110100001111000100010001110100000000000") port map( O =>C_4_S_0_L_5_out, I0 =>  inp_feat(234), I1 =>  inp_feat(464), I2 =>  inp_feat(315), I3 =>  inp_feat(71), I4 =>  inp_feat(82), I5 =>  inp_feat(74)); 
C_4_S_1_L_0_inst : LUT6 generic map(INIT => "0000010111001110110011101100000011111111111011111100111011000000") port map( O =>C_4_S_1_L_0_out, I0 =>  inp_feat(405), I1 =>  inp_feat(494), I2 =>  inp_feat(444), I3 =>  inp_feat(28), I4 =>  inp_feat(222), I5 =>  inp_feat(312)); 
C_4_S_1_L_1_inst : LUT6 generic map(INIT => "1111111001111100111111000110000011111100011011001110000010000000") port map( O =>C_4_S_1_L_1_out, I0 =>  inp_feat(153), I1 =>  inp_feat(435), I2 =>  inp_feat(71), I3 =>  inp_feat(55), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_1_L_2_inst : LUT6 generic map(INIT => "0111010111111110111111001010100001111111011010001110100000000000") port map( O =>C_4_S_1_L_2_out, I0 =>  inp_feat(234), I1 =>  inp_feat(464), I2 =>  inp_feat(315), I3 =>  inp_feat(71), I4 =>  inp_feat(74), I5 =>  inp_feat(82)); 
C_4_S_1_L_3_inst : LUT6 generic map(INIT => "1111111111101010111111100110100011101010110010001111100010000000") port map( O =>C_4_S_1_L_3_out, I0 =>  inp_feat(159), I1 =>  inp_feat(432), I2 =>  inp_feat(71), I3 =>  inp_feat(0), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_1_L_4_inst : LUT6 generic map(INIT => "1101110111111110011110101110100001111000100010001110100000000000") port map( O =>C_4_S_1_L_4_out, I0 =>  inp_feat(234), I1 =>  inp_feat(464), I2 =>  inp_feat(315), I3 =>  inp_feat(71), I4 =>  inp_feat(82), I5 =>  inp_feat(74)); 
C_4_S_1_L_5_inst : LUT6 generic map(INIT => "0111001010101000001101100010000001101000111010001010000000000000") port map( O =>C_4_S_1_L_5_out, I0 =>  inp_feat(159), I1 =>  inp_feat(436), I2 =>  inp_feat(71), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_2_L_0_inst : LUT6 generic map(INIT => "1010011011111010111111001110100001101000110010001111100010000000") port map( O =>C_4_S_2_L_0_out, I0 =>  inp_feat(159), I1 =>  inp_feat(432), I2 =>  inp_feat(71), I3 =>  inp_feat(0), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_2_L_1_inst : LUT6 generic map(INIT => "0111001111101000111111100110100011100010111010001111100010000000") port map( O =>C_4_S_2_L_1_out, I0 =>  inp_feat(159), I1 =>  inp_feat(253), I2 =>  inp_feat(71), I3 =>  inp_feat(0), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_2_L_2_inst : LUT6 generic map(INIT => "1011111000001000111110000010000001101000110010001110100000000000") port map( O =>C_4_S_2_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(432), I2 =>  inp_feat(82), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_2_L_3_inst : LUT6 generic map(INIT => "0111100001011100011110000110000011111000001011001110100010000000") port map( O =>C_4_S_2_L_3_out, I0 =>  inp_feat(153), I1 =>  inp_feat(435), I2 =>  inp_feat(71), I3 =>  inp_feat(55), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_2_L_4_inst : LUT6 generic map(INIT => "0100111011011110111011100100000001100000101010001110000000000000") port map( O =>C_4_S_2_L_4_out, I0 =>  inp_feat(432), I1 =>  inp_feat(159), I2 =>  inp_feat(82), I3 =>  inp_feat(29), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_2_L_5_inst : LUT6 generic map(INIT => "1101110100101010011111100100000011011110101010001111100000000000") port map( O =>C_4_S_2_L_5_out, I0 =>  inp_feat(15), I1 =>  inp_feat(74), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_3_L_0_inst : LUT6 generic map(INIT => "1111011010001000111110000010000001101000110010001110100000000000") port map( O =>C_4_S_3_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(432), I2 =>  inp_feat(82), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_3_L_1_inst : LUT6 generic map(INIT => "0101001100111100111111001100100001111000010000001110100010000000") port map( O =>C_4_S_3_L_1_out, I0 =>  inp_feat(52), I1 =>  inp_feat(71), I2 =>  inp_feat(385), I3 =>  inp_feat(74), I4 =>  inp_feat(170), I5 =>  inp_feat(159)); 
C_4_S_3_L_2_inst : LUT6 generic map(INIT => "1010101110110100111111001100100010111100010000001110100010000000") port map( O =>C_4_S_3_L_2_out, I0 =>  inp_feat(52), I1 =>  inp_feat(71), I2 =>  inp_feat(385), I3 =>  inp_feat(74), I4 =>  inp_feat(170), I5 =>  inp_feat(159)); 
C_4_S_3_L_3_inst : LUT6 generic map(INIT => "0011011100100100111111101010100001011111011010001110100010000000") port map( O =>C_4_S_3_L_3_out, I0 =>  inp_feat(253), I1 =>  inp_feat(0), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_3_L_4_inst : LUT6 generic map(INIT => "1011001101100110011111101010000010110111010010001110100010000000") port map( O =>C_4_S_3_L_4_out, I0 =>  inp_feat(0), I1 =>  inp_feat(435), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_3_L_5_inst : LUT6 generic map(INIT => "0110101111101100110111100000000011111111111011001110100010000000") port map( O =>C_4_S_3_L_5_out, I0 =>  inp_feat(0), I1 =>  inp_feat(15), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_4_L_0_inst : LUT6 generic map(INIT => "0000000001101000111101100010000010101000111010001010000000000000") port map( O =>C_4_S_4_L_0_out, I0 =>  inp_feat(159), I1 =>  inp_feat(436), I2 =>  inp_feat(71), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_4_L_1_inst : LUT6 generic map(INIT => "1010110111111010001111000110000001100000010010001111100010000000") port map( O =>C_4_S_4_L_1_out, I0 =>  inp_feat(159), I1 =>  inp_feat(432), I2 =>  inp_feat(71), I3 =>  inp_feat(0), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_4_L_2_inst : LUT6 generic map(INIT => "0001011001101000001110000010000010101000010010001110100000000000") port map( O =>C_4_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(432), I2 =>  inp_feat(82), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_4_L_3_inst : LUT6 generic map(INIT => "1111101011101010110010000010000001001000111010001110100000000000") port map( O =>C_4_S_4_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(432), I2 =>  inp_feat(82), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_4_L_4_inst : LUT6 generic map(INIT => "0001000101101000011111101010000000101000011010001110000000000000") port map( O =>C_4_S_4_L_4_out, I0 =>  inp_feat(159), I1 =>  inp_feat(436), I2 =>  inp_feat(71), I3 =>  inp_feat(346), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_4_L_5_inst : LUT6 generic map(INIT => "1111111110111100111111101010100011011111011010001110100010000000") port map( O =>C_4_S_4_L_5_out, I0 =>  inp_feat(253), I1 =>  inp_feat(0), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_5_L_0_inst : LUT6 generic map(INIT => "1111110110111100011111101000100001011111011010001110100010000000") port map( O =>C_4_S_5_L_0_out, I0 =>  inp_feat(253), I1 =>  inp_feat(0), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_5_L_1_inst : LUT6 generic map(INIT => "0101000000101000011111100000000001101000101010001100000010000000") port map( O =>C_4_S_5_L_1_out, I0 =>  inp_feat(15), I1 =>  inp_feat(82), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_5_L_2_inst : LUT6 generic map(INIT => "1111111100110000110111101010100011111110011010001110100010000000") port map( O =>C_4_S_5_L_2_out, I0 =>  inp_feat(253), I1 =>  inp_feat(0), I2 =>  inp_feat(153), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_5_L_3_inst : LUT6 generic map(INIT => "0111011011101000000010100010100001111000101000001011100010000000") port map( O =>C_4_S_5_L_3_out, I0 =>  inp_feat(385), I1 =>  inp_feat(170), I2 =>  inp_feat(159), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_5_L_4_inst : LUT6 generic map(INIT => "1000011000001000101000100110000010100110100011001010000000000000") port map( O =>C_4_S_5_L_4_out, I0 =>  inp_feat(159), I1 =>  inp_feat(436), I2 =>  inp_feat(346), I3 =>  inp_feat(71), I4 =>  inp_feat(52), I5 =>  inp_feat(327)); 
C_4_S_5_L_5_inst : LUT6 generic map(INIT => "0000011111100001110100001010000111111111111101111110111101000010") port map( O =>C_4_S_5_L_5_out, I0 =>  inp_feat(138), I1 =>  inp_feat(180), I2 =>  inp_feat(462), I3 =>  inp_feat(275), I4 =>  inp_feat(3), I5 =>  inp_feat(421)); 
C_5_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000000001011100000000000101110000010101111111") port map( O =>C_5_S_0_L_0_out, I0 =>  inp_feat(253), I1 =>  inp_feat(315), I2 =>  inp_feat(435), I3 =>  inp_feat(0), I4 =>  inp_feat(102), I5 =>  inp_feat(71)); 
C_5_S_0_L_1_inst : LUT6 generic map(INIT => "0000011100110010011111111110000000010111111000101111111111111001") port map( O =>C_5_S_0_L_1_out, I0 =>  inp_feat(15), I1 =>  inp_feat(325), I2 =>  inp_feat(58), I3 =>  inp_feat(497), I4 =>  inp_feat(180), I5 =>  inp_feat(29)); 
C_5_S_0_L_2_inst : LUT6 generic map(INIT => "0010111101101110101011101011111000000000001011100011011010111011") port map( O =>C_5_S_0_L_2_out, I0 =>  inp_feat(257), I1 =>  inp_feat(170), I2 =>  inp_feat(72), I3 =>  inp_feat(82), I4 =>  inp_feat(319), I5 =>  inp_feat(375)); 
C_5_S_0_L_3_inst : LUT6 generic map(INIT => "0001011100010001101101011010000001111111111111110000001010001010") port map( O =>C_5_S_0_L_3_out, I0 =>  inp_feat(410), I1 =>  inp_feat(327), I2 =>  inp_feat(234), I3 =>  inp_feat(306), I4 =>  inp_feat(320), I5 =>  inp_feat(431)); 
C_5_S_0_L_4_inst : LUT6 generic map(INIT => "0101001111110001011111111111011100000000000000000010000010101000") port map( O =>C_5_S_0_L_4_out, I0 =>  inp_feat(346), I1 =>  inp_feat(319), I2 =>  inp_feat(228), I3 =>  inp_feat(11), I4 =>  inp_feat(82), I5 =>  inp_feat(312)); 
C_5_S_0_L_5_inst : LUT6 generic map(INIT => "0100100100001011110010001100101000000000000000000000000000001000") port map( O =>C_5_S_0_L_5_out, I0 =>  inp_feat(417), I1 =>  inp_feat(177), I2 =>  inp_feat(22), I3 =>  inp_feat(254), I4 =>  inp_feat(164), I5 =>  inp_feat(312)); 
C_5_S_1_L_0_inst : LUT6 generic map(INIT => "0000011100110010011111111110000000010111111000101111111111111001") port map( O =>C_5_S_1_L_0_out, I0 =>  inp_feat(15), I1 =>  inp_feat(325), I2 =>  inp_feat(58), I3 =>  inp_feat(497), I4 =>  inp_feat(180), I5 =>  inp_feat(29)); 
C_5_S_1_L_1_inst : LUT6 generic map(INIT => "0010111101101110101011101011111000000000001011100011011010111011") port map( O =>C_5_S_1_L_1_out, I0 =>  inp_feat(257), I1 =>  inp_feat(170), I2 =>  inp_feat(72), I3 =>  inp_feat(82), I4 =>  inp_feat(319), I5 =>  inp_feat(375)); 
C_5_S_1_L_2_inst : LUT6 generic map(INIT => "0001011100010001101101011010000001111111111111110000001010001010") port map( O =>C_5_S_1_L_2_out, I0 =>  inp_feat(410), I1 =>  inp_feat(327), I2 =>  inp_feat(234), I3 =>  inp_feat(306), I4 =>  inp_feat(320), I5 =>  inp_feat(431)); 
C_5_S_1_L_3_inst : LUT6 generic map(INIT => "0101001111110001011111111111011100000000000000000010000010101000") port map( O =>C_5_S_1_L_3_out, I0 =>  inp_feat(346), I1 =>  inp_feat(319), I2 =>  inp_feat(228), I3 =>  inp_feat(11), I4 =>  inp_feat(82), I5 =>  inp_feat(312)); 
C_5_S_1_L_4_inst : LUT6 generic map(INIT => "0100100100001011110010001100101000000000000000000000000000001000") port map( O =>C_5_S_1_L_4_out, I0 =>  inp_feat(417), I1 =>  inp_feat(177), I2 =>  inp_feat(22), I3 =>  inp_feat(254), I4 =>  inp_feat(164), I5 =>  inp_feat(312)); 
C_5_S_1_L_5_inst : LUT6 generic map(INIT => "0000000110110000000000001101000011111111110000010000001010100001") port map( O =>C_5_S_1_L_5_out, I0 =>  inp_feat(139), I1 =>  inp_feat(172), I2 =>  inp_feat(204), I3 =>  inp_feat(325), I4 =>  inp_feat(58), I5 =>  inp_feat(160)); 
C_5_S_2_L_0_inst : LUT6 generic map(INIT => "0001001100011011000000000001011111111111000010010000000000000000") port map( O =>C_5_S_2_L_0_out, I0 =>  inp_feat(429), I1 =>  inp_feat(43), I2 =>  inp_feat(263), I3 =>  inp_feat(160), I4 =>  inp_feat(89), I5 =>  inp_feat(348)); 
C_5_S_2_L_1_inst : LUT6 generic map(INIT => "0011010111100001000000000010000011100101111111110000000000000000") port map( O =>C_5_S_2_L_1_out, I0 =>  inp_feat(394), I1 =>  inp_feat(71), I2 =>  inp_feat(10), I3 =>  inp_feat(410), I4 =>  inp_feat(312), I5 =>  inp_feat(92)); 
C_5_S_2_L_2_inst : LUT6 generic map(INIT => "1110111111111011000000000000010000000001000000100000000000000000") port map( O =>C_5_S_2_L_2_out, I0 =>  inp_feat(296), I1 =>  inp_feat(82), I2 =>  inp_feat(22), I3 =>  inp_feat(170), I4 =>  inp_feat(79), I5 =>  inp_feat(312)); 
C_5_S_2_L_3_inst : LUT6 generic map(INIT => "0000100000001101000011001111111111000101000111011101111111111101") port map( O =>C_5_S_2_L_3_out, I0 =>  inp_feat(0), I1 =>  inp_feat(391), I2 =>  inp_feat(82), I3 =>  inp_feat(11), I4 =>  inp_feat(253), I5 =>  inp_feat(327)); 
C_5_S_2_L_4_inst : LUT6 generic map(INIT => "0000100001010001110100000001000011010001110100010000010001110101") port map( O =>C_5_S_2_L_4_out, I0 =>  inp_feat(95), I1 =>  inp_feat(407), I2 =>  inp_feat(507), I3 =>  inp_feat(1), I4 =>  inp_feat(359), I5 =>  inp_feat(111)); 
C_5_S_2_L_5_inst : LUT6 generic map(INIT => "1101011101110011101101111111111100000000000000010000000000000111") port map( O =>C_5_S_2_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(319), I2 =>  inp_feat(0), I3 =>  inp_feat(15), I4 =>  inp_feat(410), I5 =>  inp_feat(312)); 
C_5_S_3_L_0_inst : LUT6 generic map(INIT => "0111001100010011111110110001001000000011000100100000000000000000") port map( O =>C_5_S_3_L_0_out, I0 =>  inp_feat(58), I1 =>  inp_feat(82), I2 =>  inp_feat(11), I3 =>  inp_feat(286), I4 =>  inp_feat(440), I5 =>  inp_feat(312)); 
C_5_S_3_L_1_inst : LUT6 generic map(INIT => "0000010111011001111110000000001100000000000000000000000000000000") port map( O =>C_5_S_3_L_1_out, I0 =>  inp_feat(222), I1 =>  inp_feat(310), I2 =>  inp_feat(90), I3 =>  inp_feat(410), I4 =>  inp_feat(126), I5 =>  inp_feat(312)); 
C_5_S_3_L_2_inst : LUT6 generic map(INIT => "0000010000000111010100110000110001110110000000001110101111110111") port map( O =>C_5_S_3_L_2_out, I0 =>  inp_feat(124), I1 =>  inp_feat(450), I2 =>  inp_feat(353), I3 =>  inp_feat(204), I4 =>  inp_feat(415), I5 =>  inp_feat(96)); 
C_5_S_3_L_3_inst : LUT6 generic map(INIT => "1111011110010010111111100000010000010000000000000000000000000000") port map( O =>C_5_S_3_L_3_out, I0 =>  inp_feat(71), I1 =>  inp_feat(33), I2 =>  inp_feat(389), I3 =>  inp_feat(380), I4 =>  inp_feat(23), I5 =>  inp_feat(312)); 
C_5_S_3_L_4_inst : LUT6 generic map(INIT => "1001001110001111000010110000111010111111101111110000100101010100") port map( O =>C_5_S_3_L_4_out, I0 =>  inp_feat(282), I1 =>  inp_feat(339), I2 =>  inp_feat(455), I3 =>  inp_feat(37), I4 =>  inp_feat(130), I5 =>  inp_feat(203)); 
C_5_S_3_L_5_inst : LUT6 generic map(INIT => "0010000011110000000000000001010011111001111101010101010001011000") port map( O =>C_5_S_3_L_5_out, I0 =>  inp_feat(173), I1 =>  inp_feat(233), I2 =>  inp_feat(373), I3 =>  inp_feat(29), I4 =>  inp_feat(182), I5 =>  inp_feat(403)); 
C_5_S_4_L_0_inst : LUT6 generic map(INIT => "1000100001000011000000000110010010001000100010000000000000001000") port map( O =>C_5_S_4_L_0_out, I0 =>  inp_feat(476), I1 =>  inp_feat(282), I2 =>  inp_feat(287), I3 =>  inp_feat(403), I4 =>  inp_feat(7), I5 =>  inp_feat(254)); 
C_5_S_4_L_1_inst : LUT6 generic map(INIT => "0101010101111111000110110011111100000000000100010000000000000001") port map( O =>C_5_S_4_L_1_out, I0 =>  inp_feat(180), I1 =>  inp_feat(385), I2 =>  inp_feat(164), I3 =>  inp_feat(410), I4 =>  inp_feat(254), I5 =>  inp_feat(312)); 
C_5_S_4_L_2_inst : LUT6 generic map(INIT => "1011011111011101000101110001110100000011000000000000000100000000") port map( O =>C_5_S_4_L_2_out, I0 =>  inp_feat(203), I1 =>  inp_feat(230), I2 =>  inp_feat(0), I3 =>  inp_feat(403), I4 =>  inp_feat(286), I5 =>  inp_feat(312)); 
C_5_S_4_L_3_inst : LUT6 generic map(INIT => "1000001100000111010011010000010000000001000000000001010100000000") port map( O =>C_5_S_4_L_3_out, I0 =>  inp_feat(253), I1 =>  inp_feat(124), I2 =>  inp_feat(121), I3 =>  inp_feat(38), I4 =>  inp_feat(11), I5 =>  inp_feat(391)); 
C_5_S_4_L_4_inst : LUT6 generic map(INIT => "0010000101110000011110010000000100111101000010011010110100000001") port map( O =>C_5_S_4_L_4_out, I0 =>  inp_feat(510), I1 =>  inp_feat(325), I2 =>  inp_feat(91), I3 =>  inp_feat(380), I4 =>  inp_feat(16), I5 =>  inp_feat(23)); 
C_5_S_4_L_5_inst : LUT6 generic map(INIT => "0011000110110110111001110110110100000000000000000000000000001100") port map( O =>C_5_S_4_L_5_out, I0 =>  inp_feat(249), I1 =>  inp_feat(199), I2 =>  inp_feat(71), I3 =>  inp_feat(230), I4 =>  inp_feat(0), I5 =>  inp_feat(312)); 
C_5_S_5_L_0_inst : LUT6 generic map(INIT => "0101100010011110100111011100110100000000000000000000000000001100") port map( O =>C_5_S_5_L_0_out, I0 =>  inp_feat(475), I1 =>  inp_feat(303), I2 =>  inp_feat(71), I3 =>  inp_feat(230), I4 =>  inp_feat(0), I5 =>  inp_feat(312)); 
C_5_S_5_L_1_inst : LUT6 generic map(INIT => "0010000001010001111000000100110100000000000000000000000000000000") port map( O =>C_5_S_5_L_1_out, I0 =>  inp_feat(92), I1 =>  inp_feat(387), I2 =>  inp_feat(106), I3 =>  inp_feat(301), I4 =>  inp_feat(229), I5 =>  inp_feat(312)); 
C_5_S_5_L_2_inst : LUT6 generic map(INIT => "1011111100101110001010101111111000000000000000000000000010110000") port map( O =>C_5_S_5_L_2_out, I0 =>  inp_feat(162), I1 =>  inp_feat(323), I2 =>  inp_feat(226), I3 =>  inp_feat(0), I4 =>  inp_feat(71), I5 =>  inp_feat(312)); 
C_5_S_5_L_3_inst : LUT6 generic map(INIT => "0101010000001100000010000010100011001000000000000000000000000000") port map( O =>C_5_S_5_L_3_out, I0 =>  inp_feat(58), I1 =>  inp_feat(57), I2 =>  inp_feat(353), I3 =>  inp_feat(344), I4 =>  inp_feat(342), I5 =>  inp_feat(254)); 
C_5_S_5_L_4_inst : LUT6 generic map(INIT => "1010111111101111111010111101101100000000000010010010001011111010") port map( O =>C_5_S_5_L_4_out, I0 =>  inp_feat(182), I1 =>  inp_feat(71), I2 =>  inp_feat(174), I3 =>  inp_feat(262), I4 =>  inp_feat(330), I5 =>  inp_feat(219)); 
C_5_S_5_L_5_inst : LUT6 generic map(INIT => "0101000000000000000101010001000010111101101100001111111001110111") port map( O =>C_5_S_5_L_5_out, I0 =>  inp_feat(1), I1 =>  inp_feat(113), I2 =>  inp_feat(101), I3 =>  inp_feat(510), I4 =>  inp_feat(59), I5 =>  inp_feat(242)); 
C_6_S_0_L_0_inst : LUT6 generic map(INIT => "1111110111010101111100001110000011000001010000001110100000000000") port map( O =>C_6_S_0_L_0_out, I0 =>  inp_feat(15), I1 =>  inp_feat(402), I2 =>  inp_feat(206), I3 =>  inp_feat(143), I4 =>  inp_feat(352), I5 =>  inp_feat(365)); 
C_6_S_0_L_1_inst : LUT6 generic map(INIT => "0000000011000000110011001110100011101010111011101110101011101010") port map( O =>C_6_S_0_L_1_out, I0 =>  inp_feat(222), I1 =>  inp_feat(30), I2 =>  inp_feat(274), I3 =>  inp_feat(175), I4 =>  inp_feat(230), I5 =>  inp_feat(20)); 
C_6_S_0_L_2_inst : LUT6 generic map(INIT => "1111001110110010111110100101101000110000101100001010101000101010") port map( O =>C_6_S_0_L_2_out, I0 =>  inp_feat(191), I1 =>  inp_feat(385), I2 =>  inp_feat(365), I3 =>  inp_feat(159), I4 =>  inp_feat(373), I5 =>  inp_feat(462)); 
C_6_S_0_L_3_inst : LUT6 generic map(INIT => "0001010011111101010101001011111100010000000111011100110000111111") port map( O =>C_6_S_0_L_3_out, I0 =>  inp_feat(453), I1 =>  inp_feat(397), I2 =>  inp_feat(318), I3 =>  inp_feat(289), I4 =>  inp_feat(272), I5 =>  inp_feat(454)); 
C_6_S_0_L_4_inst : LUT6 generic map(INIT => "1111110111011101000100001101010011000001000100000001000000000000") port map( O =>C_6_S_0_L_4_out, I0 =>  inp_feat(507), I1 =>  inp_feat(274), I2 =>  inp_feat(169), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_0_L_5_inst : LUT6 generic map(INIT => "1110011011101111110001001000010001001000000111110000000010000001") port map( O =>C_6_S_0_L_5_out, I0 =>  inp_feat(365), I1 =>  inp_feat(274), I2 =>  inp_feat(289), I3 =>  inp_feat(133), I4 =>  inp_feat(100), I5 =>  inp_feat(454)); 
C_6_S_1_L_0_inst : LUT6 generic map(INIT => "0000000011000000110011001110100011101010111011101110101011101010") port map( O =>C_6_S_1_L_0_out, I0 =>  inp_feat(222), I1 =>  inp_feat(30), I2 =>  inp_feat(274), I3 =>  inp_feat(175), I4 =>  inp_feat(230), I5 =>  inp_feat(20)); 
C_6_S_1_L_1_inst : LUT6 generic map(INIT => "1111001110110010111110100101101000110000101100001010101000101010") port map( O =>C_6_S_1_L_1_out, I0 =>  inp_feat(191), I1 =>  inp_feat(385), I2 =>  inp_feat(365), I3 =>  inp_feat(159), I4 =>  inp_feat(373), I5 =>  inp_feat(462)); 
C_6_S_1_L_2_inst : LUT6 generic map(INIT => "0001010011111101010101001011111100010000000111011100110000111111") port map( O =>C_6_S_1_L_2_out, I0 =>  inp_feat(453), I1 =>  inp_feat(397), I2 =>  inp_feat(318), I3 =>  inp_feat(289), I4 =>  inp_feat(272), I5 =>  inp_feat(454)); 
C_6_S_1_L_3_inst : LUT6 generic map(INIT => "1111110111011101000100001101010011000001000100000001000000000000") port map( O =>C_6_S_1_L_3_out, I0 =>  inp_feat(507), I1 =>  inp_feat(274), I2 =>  inp_feat(169), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_1_L_4_inst : LUT6 generic map(INIT => "1110011011101111110001001000010001001000000111110000000010000001") port map( O =>C_6_S_1_L_4_out, I0 =>  inp_feat(365), I1 =>  inp_feat(274), I2 =>  inp_feat(289), I3 =>  inp_feat(133), I4 =>  inp_feat(100), I5 =>  inp_feat(454)); 
C_6_S_1_L_5_inst : LUT6 generic map(INIT => "0000011011001101101011100101110100001100111101000000000011111101") port map( O =>C_6_S_1_L_5_out, I0 =>  inp_feat(144), I1 =>  inp_feat(279), I2 =>  inp_feat(70), I3 =>  inp_feat(182), I4 =>  inp_feat(277), I5 =>  inp_feat(30)); 
C_6_S_2_L_0_inst : LUT6 generic map(INIT => "1011011111110011111110011010111101110000111101001111111100110101") port map( O =>C_6_S_2_L_0_out, I0 =>  inp_feat(352), I1 =>  inp_feat(385), I2 =>  inp_feat(365), I3 =>  inp_feat(159), I4 =>  inp_feat(373), I5 =>  inp_feat(462)); 
C_6_S_2_L_1_inst : LUT6 generic map(INIT => "0010101001100110111011001110000000000000000010111111010000100000") port map( O =>C_6_S_2_L_1_out, I0 =>  inp_feat(78), I1 =>  inp_feat(365), I2 =>  inp_feat(362), I3 =>  inp_feat(70), I4 =>  inp_feat(507), I5 =>  inp_feat(30)); 
C_6_S_2_L_2_inst : LUT6 generic map(INIT => "1100111110101000101010100001000000010000101000000001000000000000") port map( O =>C_6_S_2_L_2_out, I0 =>  inp_feat(342), I1 =>  inp_feat(90), I2 =>  inp_feat(180), I3 =>  inp_feat(274), I4 =>  inp_feat(100), I5 =>  inp_feat(454)); 
C_6_S_2_L_3_inst : LUT6 generic map(INIT => "0100111111100010111100010000000001111010100000100000000000000000") port map( O =>C_6_S_2_L_3_out, I0 =>  inp_feat(262), I1 =>  inp_feat(133), I2 =>  inp_feat(274), I3 =>  inp_feat(169), I4 =>  inp_feat(423), I5 =>  inp_feat(78)); 
C_6_S_2_L_4_inst : LUT6 generic map(INIT => "1100111011001111111100111100101100110010011010100000001011111011") port map( O =>C_6_S_2_L_4_out, I0 =>  inp_feat(226), I1 =>  inp_feat(182), I2 =>  inp_feat(175), I3 =>  inp_feat(417), I4 =>  inp_feat(277), I5 =>  inp_feat(356)); 
C_6_S_2_L_5_inst : LUT6 generic map(INIT => "0000001101100100000010100010100011111011111111101111110001101000") port map( O =>C_6_S_2_L_5_out, I0 =>  inp_feat(219), I1 =>  inp_feat(187), I2 =>  inp_feat(184), I3 =>  inp_feat(224), I4 =>  inp_feat(357), I5 =>  inp_feat(456)); 
C_6_S_3_L_0_inst : LUT6 generic map(INIT => "1000011110101111000011010000101100000011110011100000100000001010") port map( O =>C_6_S_3_L_0_out, I0 =>  inp_feat(31), I1 =>  inp_feat(415), I2 =>  inp_feat(453), I3 =>  inp_feat(309), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_3_L_1_inst : LUT6 generic map(INIT => "0001111111110111001011100010101000011010011110100010001010001010") port map( O =>C_6_S_3_L_1_out, I0 =>  inp_feat(217), I1 =>  inp_feat(467), I2 =>  inp_feat(417), I3 =>  inp_feat(126), I4 =>  inp_feat(100), I5 =>  inp_feat(455)); 
C_6_S_3_L_2_inst : LUT6 generic map(INIT => "1111110101111101111110100010100001100111001011110001100000000000") port map( O =>C_6_S_3_L_2_out, I0 =>  inp_feat(444), I1 =>  inp_feat(70), I2 =>  inp_feat(480), I3 =>  inp_feat(274), I4 =>  inp_feat(100), I5 =>  inp_feat(455)); 
C_6_S_3_L_3_inst : LUT6 generic map(INIT => "0011011001110101001001101110110011111110111000001111111111111111") port map( O =>C_6_S_3_L_3_out, I0 =>  inp_feat(123), I1 =>  inp_feat(370), I2 =>  inp_feat(449), I3 =>  inp_feat(273), I4 =>  inp_feat(352), I5 =>  inp_feat(312)); 
C_6_S_3_L_4_inst : LUT6 generic map(INIT => "1100111011101000001011100000110011101000000000001000000000000000") port map( O =>C_6_S_3_L_4_out, I0 =>  inp_feat(274), I1 =>  inp_feat(100), I2 =>  inp_feat(393), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_3_L_5_inst : LUT6 generic map(INIT => "1101011000010111100111011101111000000011000100011100110110001101") port map( O =>C_6_S_3_L_5_out, I0 =>  inp_feat(257), I1 =>  inp_feat(274), I2 =>  inp_feat(91), I3 =>  inp_feat(500), I4 =>  inp_feat(99), I5 =>  inp_feat(388)); 
C_6_S_4_L_0_inst : LUT6 generic map(INIT => "1011101110110011110000101000000011101000000000000000000000000000") port map( O =>C_6_S_4_L_0_out, I0 =>  inp_feat(423), I1 =>  inp_feat(468), I2 =>  inp_feat(169), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_4_L_1_inst : LUT6 generic map(INIT => "0001001010000000010100101110001011110011000000100010000000000000") port map( O =>C_6_S_4_L_1_out, I0 =>  inp_feat(423), I1 =>  inp_feat(98), I2 =>  inp_feat(78), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_4_L_2_inst : LUT6 generic map(INIT => "1010110101010111111111110001111100001100001100000001100000000000") port map( O =>C_6_S_4_L_2_out, I0 =>  inp_feat(218), I1 =>  inp_feat(101), I2 =>  inp_feat(122), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_4_L_3_inst : LUT6 generic map(INIT => "0101100011110010110000001010000000001000110000010000000000000000") port map( O =>C_6_S_4_L_3_out, I0 =>  inp_feat(143), I1 =>  inp_feat(350), I2 =>  inp_feat(30), I3 =>  inp_feat(363), I4 =>  inp_feat(419), I5 =>  inp_feat(28)); 
C_6_S_4_L_4_inst : LUT6 generic map(INIT => "0001011100100110111101111010001011101011111100011111111111111011") port map( O =>C_6_S_4_L_4_out, I0 =>  inp_feat(203), I1 =>  inp_feat(476), I2 =>  inp_feat(28), I3 =>  inp_feat(283), I4 =>  inp_feat(157), I5 =>  inp_feat(125)); 
C_6_S_4_L_5_inst : LUT6 generic map(INIT => "1010110011110110011011100000010001011100101111110000001000000000") port map( O =>C_6_S_4_L_5_out, I0 =>  inp_feat(387), I1 =>  inp_feat(386), I2 =>  inp_feat(257), I3 =>  inp_feat(363), I4 =>  inp_feat(179), I5 =>  inp_feat(28)); 
C_6_S_5_L_0_inst : LUT6 generic map(INIT => "0011010110111111100011000010111110101101000011010010110000000000") port map( O =>C_6_S_5_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(186), I2 =>  inp_feat(182), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_5_L_1_inst : LUT6 generic map(INIT => "1101001010110001101110101010001011010010000000000011000000000000") port map( O =>C_6_S_5_L_1_out, I0 =>  inp_feat(222), I1 =>  inp_feat(380), I2 =>  inp_feat(423), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_5_L_2_inst : LUT6 generic map(INIT => "1010000010101000011000000100000000100000001011000000000010000110") port map( O =>C_6_S_5_L_2_out, I0 =>  inp_feat(194), I1 =>  inp_feat(402), I2 =>  inp_feat(301), I3 =>  inp_feat(133), I4 =>  inp_feat(180), I5 =>  inp_feat(24)); 
C_6_S_5_L_3_inst : LUT6 generic map(INIT => "0001010100111101100111100010111110101101000011010010110000000000") port map( O =>C_6_S_5_L_3_out, I0 =>  inp_feat(78), I1 =>  inp_feat(186), I2 =>  inp_feat(182), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_5_L_4_inst : LUT6 generic map(INIT => "1101101001111110001101000001110101101101000011010010110000000000") port map( O =>C_6_S_5_L_4_out, I0 =>  inp_feat(510), I1 =>  inp_feat(186), I2 =>  inp_feat(182), I3 =>  inp_feat(142), I4 =>  inp_feat(277), I5 =>  inp_feat(462)); 
C_6_S_5_L_5_inst : LUT6 generic map(INIT => "0000101111110111111111110101000101001010011110110101111101000000") port map( O =>C_6_S_5_L_5_out, I0 =>  inp_feat(485), I1 =>  inp_feat(126), I2 =>  inp_feat(173), I3 =>  inp_feat(274), I4 =>  inp_feat(423), I5 =>  inp_feat(429)); 
C_7_S_0_L_0_inst : LUT6 generic map(INIT => "1111110111010101111100001110000011000001010000001110100000000000") port map( O =>C_7_S_0_L_0_out, I0 =>  inp_feat(15), I1 =>  inp_feat(402), I2 =>  inp_feat(206), I3 =>  inp_feat(143), I4 =>  inp_feat(352), I5 =>  inp_feat(365)); 
C_7_S_0_L_1_inst : LUT6 generic map(INIT => "0101111001011111010111010100110011111111111111111101110100001111") port map( O =>C_7_S_0_L_1_out, I0 =>  inp_feat(435), I1 =>  inp_feat(262), I2 =>  inp_feat(482), I3 =>  inp_feat(28), I4 =>  inp_feat(423), I5 =>  inp_feat(183)); 
C_7_S_0_L_2_inst : LUT6 generic map(INIT => "1110111010101000101111011110000000000000100100001001011110000000") port map( O =>C_7_S_0_L_2_out, I0 =>  inp_feat(227), I1 =>  inp_feat(86), I2 =>  inp_feat(454), I3 =>  inp_feat(372), I4 =>  inp_feat(248), I5 =>  inp_feat(423)); 
C_7_S_0_L_3_inst : LUT6 generic map(INIT => "1100100010111100000000001110100000101000111010000000000011000000") port map( O =>C_7_S_0_L_3_out, I0 =>  inp_feat(78), I1 =>  inp_feat(204), I2 =>  inp_feat(423), I3 =>  inp_feat(208), I4 =>  inp_feat(28), I5 =>  inp_feat(97)); 
C_7_S_0_L_4_inst : LUT6 generic map(INIT => "0111000000101010101011010000000001010011000010000001111100000000") port map( O =>C_7_S_0_L_4_out, I0 =>  inp_feat(342), I1 =>  inp_feat(499), I2 =>  inp_feat(65), I3 =>  inp_feat(86), I4 =>  inp_feat(78), I5 =>  inp_feat(31)); 
C_7_S_0_L_5_inst : LUT6 generic map(INIT => "1100010010000111111011000001101001000110000010000000000000000000") port map( O =>C_7_S_0_L_5_out, I0 =>  inp_feat(100), I1 =>  inp_feat(499), I2 =>  inp_feat(65), I3 =>  inp_feat(31), I4 =>  inp_feat(78), I5 =>  inp_feat(86)); 
C_7_S_1_L_0_inst : LUT6 generic map(INIT => "0101111001011111010111010100110011111111111111111101110100001111") port map( O =>C_7_S_1_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(262), I2 =>  inp_feat(482), I3 =>  inp_feat(28), I4 =>  inp_feat(423), I5 =>  inp_feat(183)); 
C_7_S_1_L_1_inst : LUT6 generic map(INIT => "1110111010101000101111011110000000000000100100001001011110000000") port map( O =>C_7_S_1_L_1_out, I0 =>  inp_feat(227), I1 =>  inp_feat(86), I2 =>  inp_feat(454), I3 =>  inp_feat(372), I4 =>  inp_feat(248), I5 =>  inp_feat(423)); 
C_7_S_1_L_2_inst : LUT6 generic map(INIT => "1100100010111100000000001110100000101000111010000000000011000000") port map( O =>C_7_S_1_L_2_out, I0 =>  inp_feat(78), I1 =>  inp_feat(204), I2 =>  inp_feat(423), I3 =>  inp_feat(208), I4 =>  inp_feat(28), I5 =>  inp_feat(97)); 
C_7_S_1_L_3_inst : LUT6 generic map(INIT => "0111000000101010101011010000000001010011000010000001111100000000") port map( O =>C_7_S_1_L_3_out, I0 =>  inp_feat(342), I1 =>  inp_feat(499), I2 =>  inp_feat(65), I3 =>  inp_feat(86), I4 =>  inp_feat(78), I5 =>  inp_feat(31)); 
C_7_S_1_L_4_inst : LUT6 generic map(INIT => "1100010010000111111011000001101001000110000010000000000000000000") port map( O =>C_7_S_1_L_4_out, I0 =>  inp_feat(100), I1 =>  inp_feat(499), I2 =>  inp_feat(65), I3 =>  inp_feat(31), I4 =>  inp_feat(78), I5 =>  inp_feat(86)); 
C_7_S_1_L_5_inst : LUT6 generic map(INIT => "0011010101101100101011110000110001111111000011100000111000000000") port map( O =>C_7_S_1_L_5_out, I0 =>  inp_feat(510), I1 =>  inp_feat(365), I2 =>  inp_feat(507), I3 =>  inp_feat(78), I4 =>  inp_feat(160), I5 =>  inp_feat(100)); 
C_7_S_2_L_0_inst : LUT6 generic map(INIT => "1110111110001111111011100000111000001111000010110000111100001000") port map( O =>C_7_S_2_L_0_out, I0 =>  inp_feat(465), I1 =>  inp_feat(24), I2 =>  inp_feat(182), I3 =>  inp_feat(78), I4 =>  inp_feat(86), I5 =>  inp_feat(423)); 
C_7_S_2_L_1_inst : LUT6 generic map(INIT => "0010111010101100001000000000000000000000000000000000001000000000") port map( O =>C_7_S_2_L_1_out, I0 =>  inp_feat(86), I1 =>  inp_feat(462), I2 =>  inp_feat(498), I3 =>  inp_feat(319), I4 =>  inp_feat(423), I5 =>  inp_feat(31)); 
C_7_S_2_L_2_inst : LUT6 generic map(INIT => "0111001111010100011101110101110100010000000101101110000010000000") port map( O =>C_7_S_2_L_2_out, I0 =>  inp_feat(76), I1 =>  inp_feat(372), I2 =>  inp_feat(0), I3 =>  inp_feat(70), I4 =>  inp_feat(373), I5 =>  inp_feat(462)); 
C_7_S_2_L_3_inst : LUT6 generic map(INIT => "1110100010011100100000000000110001000010110010001000000000000000") port map( O =>C_7_S_2_L_3_out, I0 =>  inp_feat(86), I1 =>  inp_feat(342), I2 =>  inp_feat(454), I3 =>  inp_feat(373), I4 =>  inp_feat(319), I5 =>  inp_feat(462)); 
C_7_S_2_L_4_inst : LUT6 generic map(INIT => "1010100000011100111001100100010011110111110111001111111111001100") port map( O =>C_7_S_2_L_4_out, I0 =>  inp_feat(263), I1 =>  inp_feat(218), I2 =>  inp_feat(375), I3 =>  inp_feat(455), I4 =>  inp_feat(74), I5 =>  inp_feat(54)); 
C_7_S_2_L_5_inst : LUT6 generic map(INIT => "0110111000101010101011001000000000101000001010000000000000001010") port map( O =>C_7_S_2_L_5_out, I0 =>  inp_feat(86), I1 =>  inp_feat(8), I2 =>  inp_feat(348), I3 =>  inp_feat(498), I4 =>  inp_feat(423), I5 =>  inp_feat(31)); 
C_7_S_3_L_0_inst : LUT6 generic map(INIT => "1100100000000000010110000000110001000010100000001100100000000000") port map( O =>C_7_S_3_L_0_out, I0 =>  inp_feat(86), I1 =>  inp_feat(342), I2 =>  inp_feat(454), I3 =>  inp_feat(319), I4 =>  inp_feat(373), I5 =>  inp_feat(462)); 
C_7_S_3_L_1_inst : LUT6 generic map(INIT => "1001000110110011111110111110001100101110001010001010101000000000") port map( O =>C_7_S_3_L_1_out, I0 =>  inp_feat(342), I1 =>  inp_feat(54), I2 =>  inp_feat(48), I3 =>  inp_feat(319), I4 =>  inp_feat(373), I5 =>  inp_feat(462)); 
C_7_S_3_L_2_inst : LUT6 generic map(INIT => "0100000000100110011101000001110001101000000110000101000000000000") port map( O =>C_7_S_3_L_2_out, I0 =>  inp_feat(103), I1 =>  inp_feat(173), I2 =>  inp_feat(17), I3 =>  inp_feat(24), I4 =>  inp_feat(454), I5 =>  inp_feat(100)); 
C_7_S_3_L_3_inst : LUT6 generic map(INIT => "1101000011111000101010001000000010000010100010000000000010010000") port map( O =>C_7_S_3_L_3_out, I0 =>  inp_feat(342), I1 =>  inp_feat(30), I2 =>  inp_feat(86), I3 =>  inp_feat(197), I4 =>  inp_feat(454), I5 =>  inp_feat(100)); 
C_7_S_3_L_4_inst : LUT6 generic map(INIT => "0100000001011101011111101101001111101111111110111111111111111111") port map( O =>C_7_S_3_L_4_out, I0 =>  inp_feat(48), I1 =>  inp_feat(257), I2 =>  inp_feat(480), I3 =>  inp_feat(183), I4 =>  inp_feat(74), I5 =>  inp_feat(54)); 
C_7_S_3_L_5_inst : LUT6 generic map(INIT => "0001001111011011100011101100001101110111111101110000001011111111") port map( O =>C_7_S_3_L_5_out, I0 =>  inp_feat(91), I1 =>  inp_feat(182), I2 =>  inp_feat(10), I3 =>  inp_feat(366), I4 =>  inp_feat(482), I5 =>  inp_feat(101)); 
C_7_S_4_L_0_inst : LUT6 generic map(INIT => "1110111010101010101011000000110011001110000000000000100000000000") port map( O =>C_7_S_4_L_0_out, I0 =>  inp_feat(423), I1 =>  inp_feat(175), I2 =>  inp_feat(257), I3 =>  inp_feat(301), I4 =>  inp_feat(319), I5 =>  inp_feat(462)); 
C_7_S_4_L_1_inst : LUT6 generic map(INIT => "0110100011110000110100111110000000000010001100001011001100100000") port map( O =>C_7_S_4_L_1_out, I0 =>  inp_feat(97), I1 =>  inp_feat(257), I2 =>  inp_feat(454), I3 =>  inp_feat(100), I4 =>  inp_feat(112), I5 =>  inp_feat(31)); 
C_7_S_4_L_2_inst : LUT6 generic map(INIT => "1000110010001110001111110010011000010111001111110010111000100011") port map( O =>C_7_S_4_L_2_out, I0 =>  inp_feat(100), I1 =>  inp_feat(456), I2 =>  inp_feat(374), I3 =>  inp_feat(28), I4 =>  inp_feat(117), I5 =>  inp_feat(31)); 
C_7_S_4_L_3_inst : LUT6 generic map(INIT => "0010000100101001111011111100111111111110111111110100111111111111") port map( O =>C_7_S_4_L_3_out, I0 =>  inp_feat(500), I1 =>  inp_feat(456), I2 =>  inp_feat(115), I3 =>  inp_feat(307), I4 =>  inp_feat(435), I5 =>  inp_feat(417)); 
C_7_S_4_L_4_inst : LUT6 generic map(INIT => "0100100010101010011111101111110001111111111110100111111111101111") port map( O =>C_7_S_4_L_4_out, I0 =>  inp_feat(318), I1 =>  inp_feat(126), I2 =>  inp_feat(76), I3 =>  inp_feat(85), I4 =>  inp_feat(383), I5 =>  inp_feat(377)); 
C_7_S_4_L_5_inst : LUT6 generic map(INIT => "1111111010111110001111111111111100000110001111111100111111111001") port map( O =>C_7_S_4_L_5_out, I0 =>  inp_feat(375), I1 =>  inp_feat(451), I2 =>  inp_feat(199), I3 =>  inp_feat(79), I4 =>  inp_feat(492), I5 =>  inp_feat(482)); 
C_7_S_5_L_0_inst : LUT6 generic map(INIT => "1111011111010001010100100001000000100111001011011000100000000000") port map( O =>C_7_S_5_L_0_out, I0 =>  inp_feat(224), I1 =>  inp_feat(197), I2 =>  inp_feat(28), I3 =>  inp_feat(97), I4 =>  inp_feat(454), I5 =>  inp_feat(456)); 
C_7_S_5_L_1_inst : LUT6 generic map(INIT => "1001011101011110000001010011101011111110110111100101110011111100") port map( O =>C_7_S_5_L_1_out, I0 =>  inp_feat(305), I1 =>  inp_feat(95), I2 =>  inp_feat(476), I3 =>  inp_feat(139), I4 =>  inp_feat(404), I5 =>  inp_feat(87)); 
C_7_S_5_L_2_inst : LUT6 generic map(INIT => "1101010110111011011100001110100000000110111011010100000010000000") port map( O =>C_7_S_5_L_2_out, I0 =>  inp_feat(385), I1 =>  inp_feat(365), I2 =>  inp_feat(342), I3 =>  inp_feat(257), I4 =>  inp_feat(86), I5 =>  inp_feat(347)); 
C_7_S_5_L_3_inst : LUT6 generic map(INIT => "0000010000100001011111011111010111110111111101001111111100111111") port map( O =>C_7_S_5_L_3_out, I0 =>  inp_feat(260), I1 =>  inp_feat(174), I2 =>  inp_feat(76), I3 =>  inp_feat(85), I4 =>  inp_feat(377), I5 =>  inp_feat(383)); 
C_7_S_5_L_4_inst : LUT6 generic map(INIT => "0100011011111111011011111111110010011110111111101111111111111110") port map( O =>C_7_S_5_L_4_out, I0 =>  inp_feat(354), I1 =>  inp_feat(156), I2 =>  inp_feat(167), I3 =>  inp_feat(483), I4 =>  inp_feat(83), I5 =>  inp_feat(476)); 
C_7_S_5_L_5_inst : LUT6 generic map(INIT => "0100110100001101011010110101010011111110001011111111101111111111") port map( O =>C_7_S_5_L_5_out, I0 =>  inp_feat(399), I1 =>  inp_feat(29), I2 =>  inp_feat(14), I3 =>  inp_feat(25), I4 =>  inp_feat(101), I5 =>  inp_feat(83)); 
C_8_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000010011001000010001111100000111011111110111111111111111") port map( O =>C_8_S_0_L_0_out, I0 =>  inp_feat(274), I1 =>  inp_feat(86), I2 =>  inp_feat(100), I3 =>  inp_feat(206), I4 =>  inp_feat(462), I5 =>  inp_feat(365)); 
C_8_S_0_L_1_inst : LUT6 generic map(INIT => "0000011110010011100101111101011101011111101111010111111111111111") port map( O =>C_8_S_0_L_1_out, I0 =>  inp_feat(222), I1 =>  inp_feat(356), I2 =>  inp_feat(455), I3 =>  inp_feat(403), I4 =>  inp_feat(420), I5 =>  inp_feat(227)); 
C_8_S_0_L_2_inst : LUT6 generic map(INIT => "0010100100010111001001110011111100010111101111111001111110111111") port map( O =>C_8_S_0_L_2_out, I0 =>  inp_feat(30), I1 =>  inp_feat(165), I2 =>  inp_feat(423), I3 =>  inp_feat(116), I4 =>  inp_feat(55), I5 =>  inp_feat(206)); 
C_8_S_0_L_3_inst : LUT6 generic map(INIT => "0101111110111101111100100000000011111111011111111011110110110000") port map( O =>C_8_S_0_L_3_out, I0 =>  inp_feat(250), I1 =>  inp_feat(29), I2 =>  inp_feat(111), I3 =>  inp_feat(418), I4 =>  inp_feat(444), I5 =>  inp_feat(226)); 
C_8_S_0_L_4_inst : LUT6 generic map(INIT => "0100100010111011111110011111101111101001001110111111011111111111") port map( O =>C_8_S_0_L_4_out, I0 =>  inp_feat(206), I1 =>  inp_feat(423), I2 =>  inp_feat(81), I3 =>  inp_feat(178), I4 =>  inp_feat(116), I5 =>  inp_feat(176)); 
C_8_S_0_L_5_inst : LUT6 generic map(INIT => "0110011010100101110100110111111111001101000101111011111111111111") port map( O =>C_8_S_0_L_5_out, I0 =>  inp_feat(420), I1 =>  inp_feat(402), I2 =>  inp_feat(356), I3 =>  inp_feat(462), I4 =>  inp_feat(277), I5 =>  inp_feat(196)); 
C_8_S_1_L_0_inst : LUT6 generic map(INIT => "0000011110010011100101111101011101011111101111010111111111111111") port map( O =>C_8_S_1_L_0_out, I0 =>  inp_feat(222), I1 =>  inp_feat(356), I2 =>  inp_feat(455), I3 =>  inp_feat(403), I4 =>  inp_feat(420), I5 =>  inp_feat(227)); 
C_8_S_1_L_1_inst : LUT6 generic map(INIT => "0010100100010111001001110011111100010111101111111001111110111111") port map( O =>C_8_S_1_L_1_out, I0 =>  inp_feat(30), I1 =>  inp_feat(165), I2 =>  inp_feat(423), I3 =>  inp_feat(116), I4 =>  inp_feat(55), I5 =>  inp_feat(206)); 
C_8_S_1_L_2_inst : LUT6 generic map(INIT => "0101111110111101111100100000000011111111011111111011110110110000") port map( O =>C_8_S_1_L_2_out, I0 =>  inp_feat(250), I1 =>  inp_feat(29), I2 =>  inp_feat(111), I3 =>  inp_feat(418), I4 =>  inp_feat(444), I5 =>  inp_feat(226)); 
C_8_S_1_L_3_inst : LUT6 generic map(INIT => "0100100010111011111110011111101111101001001110111111011111111111") port map( O =>C_8_S_1_L_3_out, I0 =>  inp_feat(206), I1 =>  inp_feat(423), I2 =>  inp_feat(81), I3 =>  inp_feat(178), I4 =>  inp_feat(116), I5 =>  inp_feat(176)); 
C_8_S_1_L_4_inst : LUT6 generic map(INIT => "0110011010100101110100110111111111001101000101111011111111111111") port map( O =>C_8_S_1_L_4_out, I0 =>  inp_feat(420), I1 =>  inp_feat(402), I2 =>  inp_feat(356), I3 =>  inp_feat(462), I4 =>  inp_feat(277), I5 =>  inp_feat(196)); 
C_8_S_1_L_5_inst : LUT6 generic map(INIT => "0011001101011111100111110111111110111111100111111111111111111111") port map( O =>C_8_S_1_L_5_out, I0 =>  inp_feat(423), I1 =>  inp_feat(165), I2 =>  inp_feat(55), I3 =>  inp_feat(8), I4 =>  inp_feat(176), I5 =>  inp_feat(313)); 
C_8_S_2_L_0_inst : LUT6 generic map(INIT => "0010101001110111000100110111111100010011111111111011011111111111") port map( O =>C_8_S_2_L_0_out, I0 =>  inp_feat(24), I1 =>  inp_feat(423), I2 =>  inp_feat(178), I3 =>  inp_feat(116), I4 =>  inp_feat(55), I5 =>  inp_feat(206)); 
C_8_S_2_L_1_inst : LUT6 generic map(INIT => "1101010101100101111100100000000001101101011011011011001001100000") port map( O =>C_8_S_2_L_1_out, I0 =>  inp_feat(385), I1 =>  inp_feat(100), I2 =>  inp_feat(452), I3 =>  inp_feat(372), I4 =>  inp_feat(444), I5 =>  inp_feat(342)); 
C_8_S_2_L_2_inst : LUT6 generic map(INIT => "0000000100001111010011110001111110000101000101111100011101111111") port map( O =>C_8_S_2_L_2_out, I0 =>  inp_feat(274), I1 =>  inp_feat(178), I2 =>  inp_feat(116), I3 =>  inp_feat(420), I4 =>  inp_feat(144), I5 =>  inp_feat(206)); 
C_8_S_2_L_3_inst : LUT6 generic map(INIT => "0001100011111000011100011010000011011101111110011111111110111000") port map( O =>C_8_S_2_L_3_out, I0 =>  inp_feat(272), I1 =>  inp_feat(373), I2 =>  inp_feat(420), I3 =>  inp_feat(227), I4 =>  inp_feat(446), I5 =>  inp_feat(296)); 
C_8_S_2_L_4_inst : LUT6 generic map(INIT => "0100100001001000010000000000100001000100110110001111010011110000") port map( O =>C_8_S_2_L_4_out, I0 =>  inp_feat(322), I1 =>  inp_feat(276), I2 =>  inp_feat(226), I3 =>  inp_feat(440), I4 =>  inp_feat(16), I5 =>  inp_feat(468)); 
C_8_S_2_L_5_inst : LUT6 generic map(INIT => "0001000110011111011101111111111111010011110111110111011101111111") port map( O =>C_8_S_2_L_5_out, I0 =>  inp_feat(356), I1 =>  inp_feat(279), I2 =>  inp_feat(444), I3 =>  inp_feat(97), I4 =>  inp_feat(419), I5 =>  inp_feat(196)); 
C_8_S_3_L_0_inst : LUT6 generic map(INIT => "1010000111101011010100110111111101110111100111111111011101111111") port map( O =>C_8_S_3_L_0_out, I0 =>  inp_feat(128), I1 =>  inp_feat(116), I2 =>  inp_feat(423), I3 =>  inp_feat(165), I4 =>  inp_feat(55), I5 =>  inp_feat(8)); 
C_8_S_3_L_1_inst : LUT6 generic map(INIT => "0010001100000001101100111001111111100111000111011111101111111111") port map( O =>C_8_S_3_L_1_out, I0 =>  inp_feat(402), I1 =>  inp_feat(454), I2 =>  inp_feat(178), I3 =>  inp_feat(420), I4 =>  inp_feat(427), I5 =>  inp_feat(8)); 
C_8_S_3_L_2_inst : LUT6 generic map(INIT => "1011000010000011000101011111010101110010111101001111101111111111") port map( O =>C_8_S_3_L_2_out, I0 =>  inp_feat(28), I1 =>  inp_feat(205), I2 =>  inp_feat(466), I3 =>  inp_feat(165), I4 =>  inp_feat(78), I5 =>  inp_feat(55)); 
C_8_S_3_L_3_inst : LUT6 generic map(INIT => "0000000010110011001110010111011101000011111011111101111111111111") port map( O =>C_8_S_3_L_3_out, I0 =>  inp_feat(455), I1 =>  inp_feat(178), I2 =>  inp_feat(444), I3 =>  inp_feat(423), I4 =>  inp_feat(165), I5 =>  inp_feat(55)); 
C_8_S_3_L_4_inst : LUT6 generic map(INIT => "0010101011110011010101111011000001000101110100011101110100000000") port map( O =>C_8_S_3_L_4_out, I0 =>  inp_feat(81), I1 =>  inp_feat(100), I2 =>  inp_feat(151), I3 =>  inp_feat(176), I4 =>  inp_feat(210), I5 =>  inp_feat(208)); 
C_8_S_3_L_5_inst : LUT6 generic map(INIT => "0101000101010001111100110111011111101000000000101111000100110010") port map( O =>C_8_S_3_L_5_out, I0 =>  inp_feat(415), I1 =>  inp_feat(93), I2 =>  inp_feat(200), I3 =>  inp_feat(289), I4 =>  inp_feat(225), I5 =>  inp_feat(242)); 
C_8_S_4_L_0_inst : LUT6 generic map(INIT => "0001000110010011100000000000000010010101100101111000000010010000") port map( O =>C_8_S_4_L_0_out, I0 =>  inp_feat(131), I1 =>  inp_feat(65), I2 =>  inp_feat(120), I3 =>  inp_feat(372), I4 =>  inp_feat(444), I5 =>  inp_feat(342)); 
C_8_S_4_L_1_inst : LUT6 generic map(INIT => "1110111000000001111110110111011111100011000101111000011101111111") port map( O =>C_8_S_4_L_1_out, I0 =>  inp_feat(454), I1 =>  inp_feat(343), I2 =>  inp_feat(423), I3 =>  inp_feat(420), I4 =>  inp_feat(144), I5 =>  inp_feat(176)); 
C_8_S_4_L_2_inst : LUT6 generic map(INIT => "0000001011010011011001100111111111110110110111110110111111111111") port map( O =>C_8_S_4_L_2_out, I0 =>  inp_feat(96), I1 =>  inp_feat(226), I2 =>  inp_feat(402), I3 =>  inp_feat(78), I4 =>  inp_feat(204), I5 =>  inp_feat(8)); 
C_8_S_4_L_3_inst : LUT6 generic map(INIT => "0101111100000101111111011000010111110011110100101111000000000000") port map( O =>C_8_S_4_L_3_out, I0 =>  inp_feat(440), I1 =>  inp_feat(357), I2 =>  inp_feat(175), I3 =>  inp_feat(434), I4 =>  inp_feat(180), I5 =>  inp_feat(16)); 
C_8_S_4_L_4_inst : LUT6 generic map(INIT => "1001001000010001000101101001110110111111000111111101111110101111") port map( O =>C_8_S_4_L_4_out, I0 =>  inp_feat(178), I1 =>  inp_feat(454), I2 =>  inp_feat(453), I3 =>  inp_feat(42), I4 =>  inp_feat(289), I5 =>  inp_feat(210)); 
C_8_S_4_L_5_inst : LUT6 generic map(INIT => "0100001111010011100001010001011111101111011111111101111111111111") port map( O =>C_8_S_4_L_5_out, I0 =>  inp_feat(28), I1 =>  inp_feat(423), I2 =>  inp_feat(30), I3 =>  inp_feat(465), I4 =>  inp_feat(160), I5 =>  inp_feat(313)); 
C_8_S_5_L_0_inst : LUT6 generic map(INIT => "0100010001100001110100010001000110100011111110001111111100000111") port map( O =>C_8_S_5_L_0_out, I0 =>  inp_feat(342), I1 =>  inp_feat(206), I2 =>  inp_feat(97), I3 =>  inp_feat(270), I4 =>  inp_feat(444), I5 =>  inp_feat(78)); 
C_8_S_5_L_1_inst : LUT6 generic map(INIT => "0111111100101101001100100000000011111010110010000000000000000000") port map( O =>C_8_S_5_L_1_out, I0 =>  inp_feat(454), I1 =>  inp_feat(288), I2 =>  inp_feat(42), I3 =>  inp_feat(391), I4 =>  inp_feat(32), I5 =>  inp_feat(87)); 
C_8_S_5_L_2_inst : LUT6 generic map(INIT => "0101000100000000001100111111001110011101100000001011111111111111") port map( O =>C_8_S_5_L_2_out, I0 =>  inp_feat(216), I1 =>  inp_feat(463), I2 =>  inp_feat(257), I3 =>  inp_feat(163), I4 =>  inp_feat(500), I5 =>  inp_feat(476)); 
C_8_S_5_L_3_inst : LUT6 generic map(INIT => "1010000100110111101011110111010110100111100101111111111100000111") port map( O =>C_8_S_5_L_3_out, I0 =>  inp_feat(342), I1 =>  inp_feat(423), I2 =>  inp_feat(402), I3 =>  inp_feat(67), I4 =>  inp_feat(204), I5 =>  inp_feat(47)); 
C_8_S_5_L_4_inst : LUT6 generic map(INIT => "1111000100000011010000010111111110010101011111110011011111111111") port map( O =>C_8_S_5_L_4_out, I0 =>  inp_feat(274), I1 =>  inp_feat(28), I2 =>  inp_feat(444), I3 =>  inp_feat(30), I4 =>  inp_feat(277), I5 =>  inp_feat(356)); 
C_8_S_5_L_5_inst : LUT6 generic map(INIT => "0000010100110000100111110100000110110111101100111101111100000011") port map( O =>C_8_S_5_L_5_out, I0 =>  inp_feat(423), I1 =>  inp_feat(194), I2 =>  inp_feat(402), I3 =>  inp_feat(127), I4 =>  inp_feat(204), I5 =>  inp_feat(47)); 
C_9_S_0_L_0_inst : LUT6 generic map(INIT => "1111110111010101111100001110000011000001010000001110100000000000") port map( O =>C_9_S_0_L_0_out, I0 =>  inp_feat(15), I1 =>  inp_feat(402), I2 =>  inp_feat(206), I3 =>  inp_feat(143), I4 =>  inp_feat(352), I5 =>  inp_feat(365)); 
C_9_S_0_L_1_inst : LUT6 generic map(INIT => "0101000101010000111101111110101111111100111111011000111111111011") port map( O =>C_9_S_0_L_1_out, I0 =>  inp_feat(224), I1 =>  inp_feat(112), I2 =>  inp_feat(359), I3 =>  inp_feat(370), I4 =>  inp_feat(314), I5 =>  inp_feat(183)); 
C_9_S_0_L_2_inst : LUT6 generic map(INIT => "1111101001111101010101000000100011010010010100100000010100000000") port map( O =>C_9_S_0_L_2_out, I0 =>  inp_feat(22), I1 =>  inp_feat(301), I2 =>  inp_feat(204), I3 =>  inp_feat(454), I4 =>  inp_feat(342), I5 =>  inp_feat(462)); 
C_9_S_0_L_3_inst : LUT6 generic map(INIT => "0010111100001011100011000000100000101110000010110000100000000000") port map( O =>C_9_S_0_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(165), I2 =>  inp_feat(372), I3 =>  inp_feat(510), I4 =>  inp_feat(429), I5 =>  inp_feat(28)); 
C_9_S_0_L_4_inst : LUT6 generic map(INIT => "1011101110111111000110101101111100100001100111110010001000101100") port map( O =>C_9_S_0_L_4_out, I0 =>  inp_feat(189), I1 =>  inp_feat(183), I2 =>  inp_feat(249), I3 =>  inp_feat(159), I4 =>  inp_feat(429), I5 =>  inp_feat(28)); 
C_9_S_0_L_5_inst : LUT6 generic map(INIT => "0000110100001100000011000100110111101010100010101110101000000110") port map( O =>C_9_S_0_L_5_out, I0 =>  inp_feat(365), I1 =>  inp_feat(356), I2 =>  inp_feat(72), I3 =>  inp_feat(288), I4 =>  inp_feat(96), I5 =>  inp_feat(147)); 
C_9_S_1_L_0_inst : LUT6 generic map(INIT => "0101000101010000111101111110101111111100111111011000111111111011") port map( O =>C_9_S_1_L_0_out, I0 =>  inp_feat(224), I1 =>  inp_feat(112), I2 =>  inp_feat(359), I3 =>  inp_feat(370), I4 =>  inp_feat(314), I5 =>  inp_feat(183)); 
C_9_S_1_L_1_inst : LUT6 generic map(INIT => "1111101001111101010101000000100011010010010100100000010100000000") port map( O =>C_9_S_1_L_1_out, I0 =>  inp_feat(22), I1 =>  inp_feat(301), I2 =>  inp_feat(204), I3 =>  inp_feat(454), I4 =>  inp_feat(342), I5 =>  inp_feat(462)); 
C_9_S_1_L_2_inst : LUT6 generic map(INIT => "0010111100001011100011000000100000101110000010110000100000000000") port map( O =>C_9_S_1_L_2_out, I0 =>  inp_feat(100), I1 =>  inp_feat(165), I2 =>  inp_feat(372), I3 =>  inp_feat(510), I4 =>  inp_feat(429), I5 =>  inp_feat(28)); 
C_9_S_1_L_3_inst : LUT6 generic map(INIT => "1011101110111111000110101101111100100001100111110010001000101100") port map( O =>C_9_S_1_L_3_out, I0 =>  inp_feat(189), I1 =>  inp_feat(183), I2 =>  inp_feat(249), I3 =>  inp_feat(159), I4 =>  inp_feat(429), I5 =>  inp_feat(28)); 
C_9_S_1_L_4_inst : LUT6 generic map(INIT => "0000110100001100000011000100110111101010100010101110101000000110") port map( O =>C_9_S_1_L_4_out, I0 =>  inp_feat(365), I1 =>  inp_feat(356), I2 =>  inp_feat(72), I3 =>  inp_feat(288), I4 =>  inp_feat(96), I5 =>  inp_feat(147)); 
C_9_S_1_L_5_inst : LUT6 generic map(INIT => "1101010100010101000111011111010011111111111111001111110010010100") port map( O =>C_9_S_1_L_5_out, I0 =>  inp_feat(162), I1 =>  inp_feat(310), I2 =>  inp_feat(10), I3 =>  inp_feat(224), I4 =>  inp_feat(27), I5 =>  inp_feat(507)); 
C_9_S_2_L_0_inst : LUT6 generic map(INIT => "1001000111101100010001011110111100001101111110000000001010100010") port map( O =>C_9_S_2_L_0_out, I0 =>  inp_feat(303), I1 =>  inp_feat(403), I2 =>  inp_feat(369), I3 =>  inp_feat(354), I4 =>  inp_feat(100), I5 =>  inp_feat(86)); 
C_9_S_2_L_1_inst : LUT6 generic map(INIT => "1011111000111100100111000000100111010101000000000000000001000000") port map( O =>C_9_S_2_L_1_out, I0 =>  inp_feat(444), I1 =>  inp_feat(454), I2 =>  inp_feat(81), I3 =>  inp_feat(350), I4 =>  inp_feat(342), I5 =>  inp_feat(462)); 
C_9_S_2_L_2_inst : LUT6 generic map(INIT => "1101100000001000000000100000110011000011000000000000100000000000") port map( O =>C_9_S_2_L_2_out, I0 =>  inp_feat(342), I1 =>  inp_feat(59), I2 =>  inp_feat(304), I3 =>  inp_feat(189), I4 =>  inp_feat(86), I5 =>  inp_feat(347)); 
C_9_S_2_L_3_inst : LUT6 generic map(INIT => "0000111011000010110001101000010000000110000010101010011010000000") port map( O =>C_9_S_2_L_3_out, I0 =>  inp_feat(28), I1 =>  inp_feat(454), I2 =>  inp_feat(17), I3 =>  inp_feat(475), I4 =>  inp_feat(363), I5 =>  inp_feat(31)); 
C_9_S_2_L_4_inst : LUT6 generic map(INIT => "0011011110111111101000111011001100000010101000000001000000000100") port map( O =>C_9_S_2_L_4_out, I0 =>  inp_feat(274), I1 =>  inp_feat(91), I2 =>  inp_feat(350), I3 =>  inp_feat(151), I4 =>  inp_feat(10), I5 =>  inp_feat(100)); 
C_9_S_2_L_5_inst : LUT6 generic map(INIT => "1111111111011111011101101110001001110110100101110011011010110000") port map( O =>C_9_S_2_L_5_out, I0 =>  inp_feat(332), I1 =>  inp_feat(1), I2 =>  inp_feat(196), I3 =>  inp_feat(39), I4 =>  inp_feat(10), I5 =>  inp_feat(31)); 
C_9_S_3_L_0_inst : LUT6 generic map(INIT => "0101010011010100100110000000000001000101000000100001010100000000") port map( O =>C_9_S_3_L_0_out, I0 =>  inp_feat(368), I1 =>  inp_feat(262), I2 =>  inp_feat(68), I3 =>  inp_feat(10), I4 =>  inp_feat(100), I5 =>  inp_feat(86)); 
C_9_S_3_L_1_inst : LUT6 generic map(INIT => "1111100000101000000000100000110001000011000000000000100000000000") port map( O =>C_9_S_3_L_1_out, I0 =>  inp_feat(342), I1 =>  inp_feat(59), I2 =>  inp_feat(304), I3 =>  inp_feat(189), I4 =>  inp_feat(86), I5 =>  inp_feat(347)); 
C_9_S_3_L_2_inst : LUT6 generic map(INIT => "0001010100110101000100100001101110111111111110110111101110011011") port map( O =>C_9_S_3_L_2_out, I0 =>  inp_feat(171), I1 =>  inp_feat(112), I2 =>  inp_feat(52), I3 =>  inp_feat(318), I4 =>  inp_feat(288), I5 =>  inp_feat(147)); 
C_9_S_3_L_3_inst : LUT6 generic map(INIT => "0000110111111001111111011111110001100110111111111111111111111100") port map( O =>C_9_S_3_L_3_out, I0 =>  inp_feat(73), I1 =>  inp_feat(344), I2 =>  inp_feat(16), I3 =>  inp_feat(22), I4 =>  inp_feat(7), I5 =>  inp_feat(500)); 
C_9_S_3_L_4_inst : LUT6 generic map(INIT => "1110101111100000000010001001100011111110111101111110001011111000") port map( O =>C_9_S_3_L_4_out, I0 =>  inp_feat(42), I1 =>  inp_feat(356), I2 =>  inp_feat(338), I3 =>  inp_feat(140), I4 =>  inp_feat(27), I5 =>  inp_feat(507)); 
C_9_S_3_L_5_inst : LUT6 generic map(INIT => "1010000101011011101110000001101011111111111111111101101100111101") port map( O =>C_9_S_3_L_5_out, I0 =>  inp_feat(296), I1 =>  inp_feat(483), I2 =>  inp_feat(91), I3 =>  inp_feat(142), I4 =>  inp_feat(27), I5 =>  inp_feat(507)); 
C_9_S_4_L_0_inst : LUT6 generic map(INIT => "0010001001001111011000011110111110101000111111111000000011111111") port map( O =>C_9_S_4_L_0_out, I0 =>  inp_feat(100), I1 =>  inp_feat(39), I2 =>  inp_feat(116), I3 =>  inp_feat(127), I4 =>  inp_feat(5), I5 =>  inp_feat(507)); 
C_9_S_4_L_1_inst : LUT6 generic map(INIT => "1111111110100111110010111110101001011011001000010001001000000000") port map( O =>C_9_S_4_L_1_out, I0 =>  inp_feat(402), I1 =>  inp_feat(151), I2 =>  inp_feat(159), I3 =>  inp_feat(488), I4 =>  inp_feat(454), I5 =>  inp_feat(100)); 
C_9_S_4_L_2_inst : LUT6 generic map(INIT => "1000010001111000100010111010000010101001111110111111111111111111") port map( O =>C_9_S_4_L_2_out, I0 =>  inp_feat(227), I1 =>  inp_feat(157), I2 =>  inp_feat(266), I3 =>  inp_feat(318), I4 =>  inp_feat(211), I5 =>  inp_feat(14)); 
C_9_S_4_L_3_inst : LUT6 generic map(INIT => "1010010011101111001111101110111001110101000111010000001111111010") port map( O =>C_9_S_4_L_3_out, I0 =>  inp_feat(342), I1 =>  inp_feat(428), I2 =>  inp_feat(22), I3 =>  inp_feat(500), I4 =>  inp_feat(344), I5 =>  inp_feat(224)); 
C_9_S_4_L_4_inst : LUT6 generic map(INIT => "0010010101111111001001010111111111111101100010000000110011000000") port map( O =>C_9_S_4_L_4_out, I0 =>  inp_feat(149), I1 =>  inp_feat(508), I2 =>  inp_feat(346), I3 =>  inp_feat(289), I4 =>  inp_feat(133), I5 =>  inp_feat(29)); 
C_9_S_4_L_5_inst : LUT6 generic map(INIT => "1001100110011111111111011011111100001010000110111111110101000001") port map( O =>C_9_S_4_L_5_out, I0 =>  inp_feat(96), I1 =>  inp_feat(91), I2 =>  inp_feat(135), I3 =>  inp_feat(289), I4 =>  inp_feat(468), I5 =>  inp_feat(351)); 
C_9_S_5_L_0_inst : LUT6 generic map(INIT => "1001100110011111111111011011111100001010000110111111110101000001") port map( O =>C_9_S_5_L_0_out, I0 =>  inp_feat(96), I1 =>  inp_feat(91), I2 =>  inp_feat(135), I3 =>  inp_feat(289), I4 =>  inp_feat(468), I5 =>  inp_feat(351)); 
C_9_S_5_L_1_inst : LUT6 generic map(INIT => "0000001110101110110011010011110011000000111111011111111011111100") port map( O =>C_9_S_5_L_1_out, I0 =>  inp_feat(174), I1 =>  inp_feat(437), I2 =>  inp_feat(440), I3 =>  inp_feat(439), I4 =>  inp_feat(104), I5 =>  inp_feat(1)); 
C_9_S_5_L_2_inst : LUT6 generic map(INIT => "1001100100101111111111101011111000101101001011111111111101101111") port map( O =>C_9_S_5_L_2_out, I0 =>  inp_feat(100), I1 =>  inp_feat(258), I2 =>  inp_feat(468), I3 =>  inp_feat(141), I4 =>  inp_feat(20), I5 =>  inp_feat(351)); 
C_9_S_5_L_3_inst : LUT6 generic map(INIT => "1000110010100011001011011111001111110111111101111000101111111001") port map( O =>C_9_S_5_L_3_out, I0 =>  inp_feat(199), I1 =>  inp_feat(403), I2 =>  inp_feat(439), I3 =>  inp_feat(170), I4 =>  inp_feat(75), I5 =>  inp_feat(431)); 
C_9_S_5_L_4_inst : LUT6 generic map(INIT => "0101010001010111101001111111101100000100010000101101101001111111") port map( O =>C_9_S_5_L_4_out, I0 =>  inp_feat(445), I1 =>  inp_feat(112), I2 =>  inp_feat(305), I3 =>  inp_feat(139), I4 =>  inp_feat(272), I5 =>  inp_feat(95)); 
C_9_S_5_L_5_inst : LUT6 generic map(INIT => "1101110100010110110111011001111100000101000110110001111101111111") port map( O =>C_9_S_5_L_5_out, I0 =>  inp_feat(299), I1 =>  inp_feat(420), I2 =>  inp_feat(406), I3 =>  inp_feat(260), I4 =>  inp_feat(313), I5 =>  inp_feat(133)); 
C_10_S_0_L_0_inst : LUT6 generic map(INIT => "1111110111010101111100001101000011010001000000001101100000000000") port map( O =>C_10_S_0_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(402), I2 =>  inp_feat(206), I3 =>  inp_feat(143), I4 =>  inp_feat(352), I5 =>  inp_feat(365)); 
C_10_S_0_L_1_inst : LUT6 generic map(INIT => "0000110001001101000000001001010011111110110111001111000001000000") port map( O =>C_10_S_0_L_1_out, I0 =>  inp_feat(173), I1 =>  inp_feat(160), I2 =>  inp_feat(143), I3 =>  inp_feat(41), I4 =>  inp_feat(423), I5 =>  inp_feat(183)); 
C_10_S_0_L_2_inst : LUT6 generic map(INIT => "1110111011101110000000011110110000000000100001000000000010001011") port map( O =>C_10_S_0_L_2_out, I0 =>  inp_feat(222), I1 =>  inp_feat(31), I2 =>  inp_feat(437), I3 =>  inp_feat(202), I4 =>  inp_feat(160), I5 =>  inp_feat(423)); 
C_10_S_0_L_3_inst : LUT6 generic map(INIT => "0101111001010001111111110111100011111111111101011110111011111110") port map( O =>C_10_S_0_L_3_out, I0 =>  inp_feat(272), I1 =>  inp_feat(25), I2 =>  inp_feat(375), I3 =>  inp_feat(93), I4 =>  inp_feat(50), I5 =>  inp_feat(453)); 
C_10_S_0_L_4_inst : LUT6 generic map(INIT => "1100100011010100101111001110100000000010000010001111100000001000") port map( O =>C_10_S_0_L_4_out, I0 =>  inp_feat(143), I1 =>  inp_feat(342), I2 =>  inp_feat(256), I3 =>  inp_feat(358), I4 =>  inp_feat(52), I5 =>  inp_feat(28)); 
C_10_S_0_L_5_inst : LUT6 generic map(INIT => "1011000010111100111011001111100000001100011000001101110000100000") port map( O =>C_10_S_0_L_5_out, I0 =>  inp_feat(143), I1 =>  inp_feat(365), I2 =>  inp_feat(41), I3 =>  inp_feat(45), I4 =>  inp_feat(299), I5 =>  inp_feat(450)); 
C_10_S_1_L_0_inst : LUT6 generic map(INIT => "0000110001001101000000001001010011111110110111001111000001000000") port map( O =>C_10_S_1_L_0_out, I0 =>  inp_feat(173), I1 =>  inp_feat(160), I2 =>  inp_feat(143), I3 =>  inp_feat(41), I4 =>  inp_feat(423), I5 =>  inp_feat(183)); 
C_10_S_1_L_1_inst : LUT6 generic map(INIT => "1110111011101110000000011110110000000000100001000000000010001011") port map( O =>C_10_S_1_L_1_out, I0 =>  inp_feat(222), I1 =>  inp_feat(31), I2 =>  inp_feat(437), I3 =>  inp_feat(202), I4 =>  inp_feat(160), I5 =>  inp_feat(423)); 
C_10_S_1_L_2_inst : LUT6 generic map(INIT => "0101111001010001111111110111100011111111111101011110111011111110") port map( O =>C_10_S_1_L_2_out, I0 =>  inp_feat(272), I1 =>  inp_feat(25), I2 =>  inp_feat(375), I3 =>  inp_feat(93), I4 =>  inp_feat(50), I5 =>  inp_feat(453)); 
C_10_S_1_L_3_inst : LUT6 generic map(INIT => "1100100011010100101111001110100000000010000010001111100000001000") port map( O =>C_10_S_1_L_3_out, I0 =>  inp_feat(143), I1 =>  inp_feat(342), I2 =>  inp_feat(256), I3 =>  inp_feat(358), I4 =>  inp_feat(52), I5 =>  inp_feat(28)); 
C_10_S_1_L_4_inst : LUT6 generic map(INIT => "1011000010111100111011001111100000001100011000001101110000100000") port map( O =>C_10_S_1_L_4_out, I0 =>  inp_feat(143), I1 =>  inp_feat(365), I2 =>  inp_feat(41), I3 =>  inp_feat(45), I4 =>  inp_feat(299), I5 =>  inp_feat(450)); 
C_10_S_1_L_5_inst : LUT6 generic map(INIT => "0111001110010011111111110011011100010001010100001111011101010001") port map( O =>C_10_S_1_L_5_out, I0 =>  inp_feat(156), I1 =>  inp_feat(318), I2 =>  inp_feat(233), I3 =>  inp_feat(399), I4 =>  inp_feat(306), I5 =>  inp_feat(244)); 
C_10_S_2_L_0_inst : LUT6 generic map(INIT => "1100100010001100000111101111010000000000101110000110100011011110") port map( O =>C_10_S_2_L_0_out, I0 =>  inp_feat(78), I1 =>  inp_feat(423), I2 =>  inp_feat(160), I3 =>  inp_feat(282), I4 =>  inp_feat(91), I5 =>  inp_feat(454)); 
C_10_S_2_L_1_inst : LUT6 generic map(INIT => "0100010011101101101101111110001100011110001000101111001100100010") port map( O =>C_10_S_2_L_1_out, I0 =>  inp_feat(43), I1 =>  inp_feat(82), I2 =>  inp_feat(432), I3 =>  inp_feat(394), I4 =>  inp_feat(223), I5 =>  inp_feat(28)); 
C_10_S_2_L_2_inst : LUT6 generic map(INIT => "1111110101011101010001011001010001001100010100110111111100000000") port map( O =>C_10_S_2_L_2_out, I0 =>  inp_feat(386), I1 =>  inp_feat(342), I2 =>  inp_feat(202), I3 =>  inp_feat(394), I4 =>  inp_feat(223), I5 =>  inp_feat(28)); 
C_10_S_2_L_3_inst : LUT6 generic map(INIT => "0111110100111111110011110011100111111011111110110000001111111101") port map( O =>C_10_S_2_L_3_out, I0 =>  inp_feat(375), I1 =>  inp_feat(482), I2 =>  inp_feat(109), I3 =>  inp_feat(449), I4 =>  inp_feat(152), I5 =>  inp_feat(418)); 
C_10_S_2_L_4_inst : LUT6 generic map(INIT => "1111101111010111011100111011001101010101001110110011001101010001") port map( O =>C_10_S_2_L_4_out, I0 =>  inp_feat(395), I1 =>  inp_feat(354), I2 =>  inp_feat(304), I3 =>  inp_feat(202), I4 =>  inp_feat(143), I5 =>  inp_feat(189)); 
C_10_S_2_L_5_inst : LUT6 generic map(INIT => "0000001100010110000000100000101111101111011011110100001111111111") port map( O =>C_10_S_2_L_5_out, I0 =>  inp_feat(493), I1 =>  inp_feat(299), I2 =>  inp_feat(221), I3 =>  inp_feat(196), I4 =>  inp_feat(388), I5 =>  inp_feat(453)); 
C_10_S_3_L_0_inst : LUT6 generic map(INIT => "0010000110010001000111011101000111110011111100111111111101010000") port map( O =>C_10_S_3_L_0_out, I0 =>  inp_feat(432), I1 =>  inp_feat(102), I2 =>  inp_feat(28), I3 =>  inp_feat(144), I4 =>  inp_feat(449), I5 =>  inp_feat(451)); 
C_10_S_3_L_1_inst : LUT6 generic map(INIT => "1100010110110111111111011111111101000101101100001101001011101010") port map( O =>C_10_S_3_L_1_out, I0 =>  inp_feat(416), I1 =>  inp_feat(76), I2 =>  inp_feat(160), I3 =>  inp_feat(52), I4 =>  inp_feat(91), I5 =>  inp_feat(429)); 
C_10_S_3_L_2_inst : LUT6 generic map(INIT => "0001000110100111011100111111111111110111001111111101111111111111") port map( O =>C_10_S_3_L_2_out, I0 =>  inp_feat(73), I1 =>  inp_feat(481), I2 =>  inp_feat(433), I3 =>  inp_feat(212), I4 =>  inp_feat(16), I5 =>  inp_feat(192)); 
C_10_S_3_L_3_inst : LUT6 generic map(INIT => "1100010111111001111111101111110000000011001010111111101011111011") port map( O =>C_10_S_3_L_3_out, I0 =>  inp_feat(476), I1 =>  inp_feat(403), I2 =>  inp_feat(300), I3 =>  inp_feat(334), I4 =>  inp_feat(188), I5 =>  inp_feat(34)); 
C_10_S_3_L_4_inst : LUT6 generic map(INIT => "1100100011101110111110111110100000000000000010001100100100100000") port map( O =>C_10_S_3_L_4_out, I0 =>  inp_feat(420), I1 =>  inp_feat(28), I2 =>  inp_feat(465), I3 =>  inp_feat(156), I4 =>  inp_feat(223), I5 =>  inp_feat(189)); 
C_10_S_3_L_5_inst : LUT6 generic map(INIT => "0001011000000011001101010000111100011001111011111111111011111111") port map( O =>C_10_S_3_L_5_out, I0 =>  inp_feat(480), I1 =>  inp_feat(43), I2 =>  inp_feat(453), I3 =>  inp_feat(257), I4 =>  inp_feat(48), I5 =>  inp_feat(269)); 
C_10_S_4_L_0_inst : LUT6 generic map(INIT => "0101011011011111010111011101111111011111011111011100100000000000") port map( O =>C_10_S_4_L_0_out, I0 =>  inp_feat(50), I1 =>  inp_feat(222), I2 =>  inp_feat(18), I3 =>  inp_feat(175), I4 =>  inp_feat(94), I5 =>  inp_feat(276)); 
C_10_S_4_L_1_inst : LUT6 generic map(INIT => "0100101111111100001011010110111111101111111111000010101111111010") port map( O =>C_10_S_4_L_1_out, I0 =>  inp_feat(378), I1 =>  inp_feat(288), I2 =>  inp_feat(67), I3 =>  inp_feat(164), I4 =>  inp_feat(71), I5 =>  inp_feat(306)); 
C_10_S_4_L_2_inst : LUT6 generic map(INIT => "1001101110111010010111011011111010111011101111110010100000000001") port map( O =>C_10_S_4_L_2_out, I0 =>  inp_feat(352), I1 =>  inp_feat(126), I2 =>  inp_feat(417), I3 =>  inp_feat(203), I4 =>  inp_feat(129), I5 =>  inp_feat(125)); 
C_10_S_4_L_3_inst : LUT6 generic map(INIT => "0010000001011011000011000001011110101101101110111001010010001011") port map( O =>C_10_S_4_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(226), I2 =>  inp_feat(306), I3 =>  inp_feat(126), I4 =>  inp_feat(456), I5 =>  inp_feat(173)); 
C_10_S_4_L_4_inst : LUT6 generic map(INIT => "1010001010110010111111001100101011101110111111101111111110111110") port map( O =>C_10_S_4_L_4_out, I0 =>  inp_feat(72), I1 =>  inp_feat(45), I2 =>  inp_feat(408), I3 =>  inp_feat(128), I4 =>  inp_feat(407), I5 =>  inp_feat(125)); 
C_10_S_4_L_5_inst : LUT6 generic map(INIT => "0000111100011100011011110011010111101110110101001111111101111111") port map( O =>C_10_S_4_L_5_out, I0 =>  inp_feat(214), I1 =>  inp_feat(406), I2 =>  inp_feat(308), I3 =>  inp_feat(128), I4 =>  inp_feat(407), I5 =>  inp_feat(125)); 
C_10_S_5_L_0_inst : LUT6 generic map(INIT => "1111101111101110010111111111111101000001010101100000111011111101") port map( O =>C_10_S_5_L_0_out, I0 =>  inp_feat(359), I1 =>  inp_feat(389), I2 =>  inp_feat(453), I3 =>  inp_feat(181), I4 =>  inp_feat(299), I5 =>  inp_feat(388)); 
C_10_S_5_L_1_inst : LUT6 generic map(INIT => "0010011011101100000100100100100011101111100010000000110010011000") port map( O =>C_10_S_5_L_1_out, I0 =>  inp_feat(78), I1 =>  inp_feat(116), I2 =>  inp_feat(449), I3 =>  inp_feat(64), I4 =>  inp_feat(256), I5 =>  inp_feat(506)); 
C_10_S_5_L_2_inst : LUT6 generic map(INIT => "0011000100111110110010101110110011011101001011101110110011011000") port map( O =>C_10_S_5_L_2_out, I0 =>  inp_feat(143), I1 =>  inp_feat(70), I2 =>  inp_feat(208), I3 =>  inp_feat(157), I4 =>  inp_feat(221), I5 =>  inp_feat(299)); 
C_10_S_5_L_3_inst : LUT6 generic map(INIT => "1111111011111111010011110101111100111100111111010100111001000100") port map( O =>C_10_S_5_L_3_out, I0 =>  inp_feat(322), I1 =>  inp_feat(195), I2 =>  inp_feat(507), I3 =>  inp_feat(224), I4 =>  inp_feat(496), I5 =>  inp_feat(247)); 
C_10_S_5_L_4_inst : LUT6 generic map(INIT => "0000001100011001110101011111100011111011111110101111000000010000") port map( O =>C_10_S_5_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(93), I2 =>  inp_feat(95), I3 =>  inp_feat(374), I4 =>  inp_feat(402), I5 =>  inp_feat(188)); 
C_10_S_5_L_5_inst : LUT6 generic map(INIT => "1101101110010111011011101111101001010001110100010100110011001100") port map( O =>C_10_S_5_L_5_out, I0 =>  inp_feat(190), I1 =>  inp_feat(330), I2 =>  inp_feat(72), I3 =>  inp_feat(399), I4 =>  inp_feat(58), I5 =>  inp_feat(86)); 
C_11_S_0_L_0_inst : LUT6 generic map(INIT => "1111110111010101111100001110000011000001010000001110100000000000") port map( O =>C_11_S_0_L_0_out, I0 =>  inp_feat(15), I1 =>  inp_feat(402), I2 =>  inp_feat(206), I3 =>  inp_feat(143), I4 =>  inp_feat(352), I5 =>  inp_feat(365)); 
C_11_S_0_L_1_inst : LUT6 generic map(INIT => "1110000011000000011011001110010000000000100000000001100011110100") port map( O =>C_11_S_0_L_1_out, I0 =>  inp_feat(454), I1 =>  inp_feat(165), I2 =>  inp_feat(423), I3 =>  inp_feat(371), I4 =>  inp_feat(91), I5 =>  inp_feat(274)); 
C_11_S_0_L_2_inst : LUT6 generic map(INIT => "1111110111000110111111110101111000011100010001001111111011011011") port map( O =>C_11_S_0_L_2_out, I0 =>  inp_feat(460), I1 =>  inp_feat(126), I2 =>  inp_feat(115), I3 =>  inp_feat(43), I4 =>  inp_feat(273), I5 =>  inp_feat(160)); 
C_11_S_0_L_3_inst : LUT6 generic map(INIT => "0110010011010100110111001101111111111111111111000111111111111111") port map( O =>C_11_S_0_L_3_out, I0 =>  inp_feat(449), I1 =>  inp_feat(318), I2 =>  inp_feat(168), I3 =>  inp_feat(322), I4 =>  inp_feat(228), I5 =>  inp_feat(183)); 
C_11_S_0_L_4_inst : LUT6 generic map(INIT => "1001001101001100111111101110100011011111010111111011000000000000") port map( O =>C_11_S_0_L_4_out, I0 =>  inp_feat(105), I1 =>  inp_feat(78), I2 =>  inp_feat(290), I3 =>  inp_feat(423), I4 =>  inp_feat(402), I5 =>  inp_feat(91)); 
C_11_S_0_L_5_inst : LUT6 generic map(INIT => "0011011010100111101111111111010011111111111101011111100101110011") port map( O =>C_11_S_0_L_5_out, I0 =>  inp_feat(361), I1 =>  inp_feat(398), I2 =>  inp_feat(142), I3 =>  inp_feat(258), I4 =>  inp_feat(329), I5 =>  inp_feat(323)); 
C_11_S_1_L_0_inst : LUT6 generic map(INIT => "1110000011000000011011001110010000000000100000000001100011110100") port map( O =>C_11_S_1_L_0_out, I0 =>  inp_feat(454), I1 =>  inp_feat(165), I2 =>  inp_feat(423), I3 =>  inp_feat(371), I4 =>  inp_feat(91), I5 =>  inp_feat(274)); 
C_11_S_1_L_1_inst : LUT6 generic map(INIT => "1111110111000110111111110101111000011100010001001111111011011011") port map( O =>C_11_S_1_L_1_out, I0 =>  inp_feat(460), I1 =>  inp_feat(126), I2 =>  inp_feat(115), I3 =>  inp_feat(43), I4 =>  inp_feat(273), I5 =>  inp_feat(160)); 
C_11_S_1_L_2_inst : LUT6 generic map(INIT => "0110010011010100110111001101111111111111111111000111111111111111") port map( O =>C_11_S_1_L_2_out, I0 =>  inp_feat(449), I1 =>  inp_feat(318), I2 =>  inp_feat(168), I3 =>  inp_feat(322), I4 =>  inp_feat(228), I5 =>  inp_feat(183)); 
C_11_S_1_L_3_inst : LUT6 generic map(INIT => "1001001101001100111111101110100011011111010111111011000000000000") port map( O =>C_11_S_1_L_3_out, I0 =>  inp_feat(105), I1 =>  inp_feat(78), I2 =>  inp_feat(290), I3 =>  inp_feat(423), I4 =>  inp_feat(402), I5 =>  inp_feat(91)); 
C_11_S_1_L_4_inst : LUT6 generic map(INIT => "0011011010100111101111111111010011111111111101011111100101110011") port map( O =>C_11_S_1_L_4_out, I0 =>  inp_feat(361), I1 =>  inp_feat(398), I2 =>  inp_feat(142), I3 =>  inp_feat(258), I4 =>  inp_feat(329), I5 =>  inp_feat(323)); 
C_11_S_1_L_5_inst : LUT6 generic map(INIT => "1100111011111011111111111111101100111101110111001111110111111101") port map( O =>C_11_S_1_L_5_out, I0 =>  inp_feat(339), I1 =>  inp_feat(486), I2 =>  inp_feat(131), I3 =>  inp_feat(200), I4 =>  inp_feat(85), I5 =>  inp_feat(357)); 
C_11_S_2_L_0_inst : LUT6 generic map(INIT => "1111110011111101111011111111001000010100111001001111111110011100") port map( O =>C_11_S_2_L_0_out, I0 =>  inp_feat(114), I1 =>  inp_feat(244), I2 =>  inp_feat(328), I3 =>  inp_feat(190), I4 =>  inp_feat(273), I5 =>  inp_feat(429)); 
C_11_S_2_L_1_inst : LUT6 generic map(INIT => "0000000110101010001011111111101110111101111111111111101101001011") port map( O =>C_11_S_2_L_1_out, I0 =>  inp_feat(288), I1 =>  inp_feat(65), I2 =>  inp_feat(174), I3 =>  inp_feat(228), I4 =>  inp_feat(511), I5 =>  inp_feat(89)); 
C_11_S_2_L_2_inst : LUT6 generic map(INIT => "1010000010111101010001001111011110011000101010101011011110100010") port map( O =>C_11_S_2_L_2_out, I0 =>  inp_feat(231), I1 =>  inp_feat(169), I2 =>  inp_feat(343), I3 =>  inp_feat(354), I4 =>  inp_feat(78), I5 =>  inp_feat(402)); 
C_11_S_2_L_3_inst : LUT6 generic map(INIT => "1010101011110010000111010111111010011111111111111101100011101111") port map( O =>C_11_S_2_L_3_out, I0 =>  inp_feat(454), I1 =>  inp_feat(442), I2 =>  inp_feat(24), I3 =>  inp_feat(393), I4 =>  inp_feat(497), I5 =>  inp_feat(91)); 
C_11_S_2_L_4_inst : LUT6 generic map(INIT => "0100010101011010000010101010001011011000111000000000000011000000") port map( O =>C_11_S_2_L_4_out, I0 =>  inp_feat(365), I1 =>  inp_feat(342), I2 =>  inp_feat(424), I3 =>  inp_feat(230), I4 =>  inp_feat(58), I5 =>  inp_feat(402)); 
C_11_S_2_L_5_inst : LUT6 generic map(INIT => "0000011110100110111110100010111111101101101111111111110111111101") port map( O =>C_11_S_2_L_5_out, I0 =>  inp_feat(174), I1 =>  inp_feat(391), I2 =>  inp_feat(16), I3 =>  inp_feat(120), I4 =>  inp_feat(290), I5 =>  inp_feat(389)); 
C_11_S_3_L_0_inst : LUT6 generic map(INIT => "1101111100111111111111111111010100111101110111100110011111010001") port map( O =>C_11_S_3_L_0_out, I0 =>  inp_feat(17), I1 =>  inp_feat(135), I2 =>  inp_feat(199), I3 =>  inp_feat(466), I4 =>  inp_feat(367), I5 =>  inp_feat(357)); 
C_11_S_3_L_1_inst : LUT6 generic map(INIT => "0000101111101011001011011111100011111111111100100110110111110111") port map( O =>C_11_S_3_L_1_out, I0 =>  inp_feat(106), I1 =>  inp_feat(128), I2 =>  inp_feat(131), I3 =>  inp_feat(200), I4 =>  inp_feat(43), I5 =>  inp_feat(273)); 
C_11_S_3_L_2_inst : LUT6 generic map(INIT => "0010110101111111111101111111111011111111010011011111110111111111") port map( O =>C_11_S_3_L_2_out, I0 =>  inp_feat(123), I1 =>  inp_feat(394), I2 =>  inp_feat(387), I3 =>  inp_feat(75), I4 =>  inp_feat(311), I5 =>  inp_feat(413)); 
C_11_S_3_L_3_inst : LUT6 generic map(INIT => "1111011100011011111011111111110011111110101010101111111110101010") port map( O =>C_11_S_3_L_3_out, I0 =>  inp_feat(511), I1 =>  inp_feat(435), I2 =>  inp_feat(62), I3 =>  inp_feat(12), I4 =>  inp_feat(107), I5 =>  inp_feat(389)); 
C_11_S_3_L_4_inst : LUT6 generic map(INIT => "0000111100001011110011011111001010111011000100111111101111111111") port map( O =>C_11_S_3_L_4_out, I0 =>  inp_feat(342), I1 =>  inp_feat(177), I2 =>  inp_feat(313), I3 =>  inp_feat(142), I4 =>  inp_feat(50), I5 =>  inp_feat(202)); 
C_11_S_3_L_5_inst : LUT6 generic map(INIT => "1110111110011100111111100000100000010110000010000010111110110000") port map( O =>C_11_S_3_L_5_out, I0 =>  inp_feat(92), I1 =>  inp_feat(402), I2 =>  inp_feat(287), I3 =>  inp_feat(342), I4 =>  inp_feat(275), I5 =>  inp_feat(100)); 
C_11_S_4_L_0_inst : LUT6 generic map(INIT => "0010000000101010000000001110100111111110111011101111011010101100") port map( O =>C_11_S_4_L_0_out, I0 =>  inp_feat(343), I1 =>  inp_feat(30), I2 =>  inp_feat(288), I3 =>  inp_feat(195), I4 =>  inp_feat(511), I5 =>  inp_feat(89)); 
C_11_S_4_L_1_inst : LUT6 generic map(INIT => "0001110110110101111111110111110111011101100111111111111111111010") port map( O =>C_11_S_4_L_1_out, I0 =>  inp_feat(445), I1 =>  inp_feat(106), I2 =>  inp_feat(45), I3 =>  inp_feat(357), I4 =>  inp_feat(138), I5 =>  inp_feat(81)); 
C_11_S_4_L_2_inst : LUT6 generic map(INIT => "1111110010001110001111101000111111101111111111111111111111000110") port map( O =>C_11_S_4_L_2_out, I0 =>  inp_feat(174), I1 =>  inp_feat(120), I2 =>  inp_feat(226), I3 =>  inp_feat(173), I4 =>  inp_feat(409), I5 =>  inp_feat(413)); 
C_11_S_4_L_3_inst : LUT6 generic map(INIT => "0110001110011111001001011111001111101101110111101000100111111111") port map( O =>C_11_S_4_L_3_out, I0 =>  inp_feat(339), I1 =>  inp_feat(120), I2 =>  inp_feat(446), I3 =>  inp_feat(344), I4 =>  inp_feat(133), I5 =>  inp_feat(393)); 
C_11_S_4_L_4_inst : LUT6 generic map(INIT => "1101011110111100101111111111100011111110111110000110111011111100") port map( O =>C_11_S_4_L_4_out, I0 =>  inp_feat(22), I1 =>  inp_feat(8), I2 =>  inp_feat(339), I3 =>  inp_feat(436), I4 =>  inp_feat(242), I5 =>  inp_feat(323)); 
C_11_S_4_L_5_inst : LUT6 generic map(INIT => "0110011101110111011101011111111011111111111111110110111111111111") port map( O =>C_11_S_4_L_5_out, I0 =>  inp_feat(413), I1 =>  inp_feat(167), I2 =>  inp_feat(248), I3 =>  inp_feat(127), I4 =>  inp_feat(94), I5 =>  inp_feat(249)); 
C_11_S_5_L_0_inst : LUT6 generic map(INIT => "1110111010101011000001001101000111111010111011101111001010000000") port map( O =>C_11_S_5_L_0_out, I0 =>  inp_feat(462), I1 =>  inp_feat(209), I2 =>  inp_feat(420), I3 =>  inp_feat(165), I4 =>  inp_feat(394), I5 =>  inp_feat(506)); 
C_11_S_5_L_1_inst : LUT6 generic map(INIT => "0011011100011010101011011001100011101000100110001100100001000100") port map( O =>C_11_S_5_L_1_out, I0 =>  inp_feat(429), I1 =>  inp_feat(365), I2 =>  inp_feat(99), I3 =>  inp_feat(165), I4 =>  inp_feat(394), I5 =>  inp_feat(506)); 
C_11_S_5_L_2_inst : LUT6 generic map(INIT => "1001111010101110110111111001100111111111110111111111100111101111") port map( O =>C_11_S_5_L_2_out, I0 =>  inp_feat(43), I1 =>  inp_feat(37), I2 =>  inp_feat(322), I3 =>  inp_feat(214), I4 =>  inp_feat(168), I5 =>  inp_feat(436)); 
C_11_S_5_L_3_inst : LUT6 generic map(INIT => "0000001111111000110011100001111111111111111100100110111111110000") port map( O =>C_11_S_5_L_3_out, I0 =>  inp_feat(26), I1 =>  inp_feat(199), I2 =>  inp_feat(330), I3 =>  inp_feat(214), I4 =>  inp_feat(318), I5 =>  inp_feat(436)); 
C_11_S_5_L_4_inst : LUT6 generic map(INIT => "1110001101011000111000001000101111111011110000001101111011000000") port map( O =>C_11_S_5_L_4_out, I0 =>  inp_feat(455), I1 =>  inp_feat(454), I2 =>  inp_feat(31), I3 =>  inp_feat(296), I4 =>  inp_feat(394), I5 =>  inp_feat(345)); 
C_11_S_5_L_5_inst : LUT6 generic map(INIT => "0100001111010100111101010000000011101010110000001100100011000000") port map( O =>C_11_S_5_L_5_out, I0 =>  inp_feat(206), I1 =>  inp_feat(342), I2 =>  inp_feat(423), I3 =>  inp_feat(408), I4 =>  inp_feat(394), I5 =>  inp_feat(345)); 
C_12_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000010000000110001111100000100011111110111111111111111") port map( O =>C_12_S_0_L_0_out, I0 =>  inp_feat(485), I1 =>  inp_feat(306), I2 =>  inp_feat(392), I3 =>  inp_feat(108), I4 =>  inp_feat(248), I5 =>  inp_feat(239)); 
C_12_S_0_L_1_inst : LUT6 generic map(INIT => "0001000000001101001111111100111110101000110010001111000000111010") port map( O =>C_12_S_0_L_1_out, I0 =>  inp_feat(304), I1 =>  inp_feat(393), I2 =>  inp_feat(288), I3 =>  inp_feat(350), I4 =>  inp_feat(194), I5 =>  inp_feat(497)); 
C_12_S_0_L_2_inst : LUT6 generic map(INIT => "0101110001111101011011111111110111111101111011011101111111011111") port map( O =>C_12_S_0_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(78), I2 =>  inp_feat(215), I3 =>  inp_feat(510), I4 =>  inp_feat(186), I5 =>  inp_feat(403)); 
C_12_S_0_L_3_inst : LUT6 generic map(INIT => "1011110011111100010011001110111010100100111111110100110111011101") port map( O =>C_12_S_0_L_3_out, I0 =>  inp_feat(239), I1 =>  inp_feat(289), I2 =>  inp_feat(186), I3 =>  inp_feat(445), I4 =>  inp_feat(149), I5 =>  inp_feat(485)); 
C_12_S_0_L_4_inst : LUT6 generic map(INIT => "0000100010011001100000001111110110111100100111100000110011101110") port map( O =>C_12_S_0_L_4_out, I0 =>  inp_feat(292), I1 =>  inp_feat(21), I2 =>  inp_feat(392), I3 =>  inp_feat(186), I4 =>  inp_feat(149), I5 =>  inp_feat(485)); 
C_12_S_0_L_5_inst : LUT6 generic map(INIT => "1001010100000100011110011111101110110000001000011110001111111111") port map( O =>C_12_S_0_L_5_out, I0 =>  inp_feat(331), I1 =>  inp_feat(123), I2 =>  inp_feat(423), I3 =>  inp_feat(186), I4 =>  inp_feat(215), I5 =>  inp_feat(211)); 
C_12_S_1_L_0_inst : LUT6 generic map(INIT => "0001000000001101001111111100111110101000110010001111000000111010") port map( O =>C_12_S_1_L_0_out, I0 =>  inp_feat(304), I1 =>  inp_feat(393), I2 =>  inp_feat(288), I3 =>  inp_feat(350), I4 =>  inp_feat(194), I5 =>  inp_feat(497)); 
C_12_S_1_L_1_inst : LUT6 generic map(INIT => "0101110001111101011011111111110111111101111011011101111111011111") port map( O =>C_12_S_1_L_1_out, I0 =>  inp_feat(190), I1 =>  inp_feat(78), I2 =>  inp_feat(215), I3 =>  inp_feat(510), I4 =>  inp_feat(186), I5 =>  inp_feat(403)); 
C_12_S_1_L_2_inst : LUT6 generic map(INIT => "1011110011111100010011001110111010100100111111110100110111011101") port map( O =>C_12_S_1_L_2_out, I0 =>  inp_feat(239), I1 =>  inp_feat(289), I2 =>  inp_feat(186), I3 =>  inp_feat(445), I4 =>  inp_feat(149), I5 =>  inp_feat(485)); 
C_12_S_1_L_3_inst : LUT6 generic map(INIT => "0000100010011001100000001111110110111100100111100000110011101110") port map( O =>C_12_S_1_L_3_out, I0 =>  inp_feat(292), I1 =>  inp_feat(21), I2 =>  inp_feat(392), I3 =>  inp_feat(186), I4 =>  inp_feat(149), I5 =>  inp_feat(485)); 
C_12_S_1_L_4_inst : LUT6 generic map(INIT => "1001010100000100011110011111101110110000001000011110001111111111") port map( O =>C_12_S_1_L_4_out, I0 =>  inp_feat(331), I1 =>  inp_feat(123), I2 =>  inp_feat(423), I3 =>  inp_feat(186), I4 =>  inp_feat(215), I5 =>  inp_feat(211)); 
C_12_S_1_L_5_inst : LUT6 generic map(INIT => "0101110111010100110001000100011111101100000000011110110010000000") port map( O =>C_12_S_1_L_5_out, I0 =>  inp_feat(168), I1 =>  inp_feat(51), I2 =>  inp_feat(257), I3 =>  inp_feat(289), I4 =>  inp_feat(215), I5 =>  inp_feat(241)); 
C_12_S_2_L_0_inst : LUT6 generic map(INIT => "1001000111110001111100001111001011111100111100001111001011110100") port map( O =>C_12_S_2_L_0_out, I0 =>  inp_feat(282), I1 =>  inp_feat(417), I2 =>  inp_feat(312), I3 =>  inp_feat(431), I4 =>  inp_feat(352), I5 =>  inp_feat(353)); 
C_12_S_2_L_1_inst : LUT6 generic map(INIT => "0101000000010101110110010000000010011000000000001100110011000000") port map( O =>C_12_S_2_L_1_out, I0 =>  inp_feat(346), I1 =>  inp_feat(451), I2 =>  inp_feat(257), I3 =>  inp_feat(276), I4 =>  inp_feat(215), I5 =>  inp_feat(211)); 
C_12_S_2_L_2_inst : LUT6 generic map(INIT => "1000001110010111000101111111011111011101110111110011111111111111") port map( O =>C_12_S_2_L_2_out, I0 =>  inp_feat(215), I1 =>  inp_feat(431), I2 =>  inp_feat(393), I3 =>  inp_feat(445), I4 =>  inp_feat(149), I5 =>  inp_feat(103)); 
C_12_S_2_L_3_inst : LUT6 generic map(INIT => "0000110100100000011000101110000001100110101000001011000010110010") port map( O =>C_12_S_2_L_3_out, I0 =>  inp_feat(289), I1 =>  inp_feat(321), I2 =>  inp_feat(296), I3 =>  inp_feat(186), I4 =>  inp_feat(215), I5 =>  inp_feat(393)); 
C_12_S_2_L_4_inst : LUT6 generic map(INIT => "1001010100011101011111011111111111101100110111010001111101111111") port map( O =>C_12_S_2_L_4_out, I0 =>  inp_feat(403), I1 =>  inp_feat(248), I2 =>  inp_feat(239), I3 =>  inp_feat(186), I4 =>  inp_feat(149), I5 =>  inp_feat(485)); 
C_12_S_2_L_5_inst : LUT6 generic map(INIT => "1000101010001000100011101000100000010000000000000000101000000000") port map( O =>C_12_S_2_L_5_out, I0 =>  inp_feat(322), I1 =>  inp_feat(131), I2 =>  inp_feat(497), I3 =>  inp_feat(149), I4 =>  inp_feat(485), I5 =>  inp_feat(73)); 
C_12_S_3_L_0_inst : LUT6 generic map(INIT => "0101010111000010001010111010000010110001111100001110100011100000") port map( O =>C_12_S_3_L_0_out, I0 =>  inp_feat(178), I1 =>  inp_feat(105), I2 =>  inp_feat(499), I3 =>  inp_feat(190), I4 =>  inp_feat(279), I5 =>  inp_feat(352)); 
C_12_S_3_L_1_inst : LUT6 generic map(INIT => "0011000001010000011110000111000110110000111100010111000011110101") port map( O =>C_12_S_3_L_1_out, I0 =>  inp_feat(334), I1 =>  inp_feat(403), I2 =>  inp_feat(312), I3 =>  inp_feat(211), I4 =>  inp_feat(279), I5 =>  inp_feat(445)); 
C_12_S_3_L_2_inst : LUT6 generic map(INIT => "1101101001101000001100101111101111011000111110111111101011111111") port map( O =>C_12_S_3_L_2_out, I0 =>  inp_feat(318), I1 =>  inp_feat(392), I2 =>  inp_feat(383), I3 =>  inp_feat(215), I4 =>  inp_feat(186), I5 =>  inp_feat(29)); 
C_12_S_3_L_3_inst : LUT6 generic map(INIT => "1000010100000111010001110001111101000111011101111111111111111111") port map( O =>C_12_S_3_L_3_out, I0 =>  inp_feat(353), I1 =>  inp_feat(306), I2 =>  inp_feat(431), I3 =>  inp_feat(510), I4 =>  inp_feat(215), I5 =>  inp_feat(186)); 
C_12_S_3_L_4_inst : LUT6 generic map(INIT => "0010000000001010101011100001001011001110000000101010101100001010") port map( O =>C_12_S_3_L_4_out, I0 =>  inp_feat(453), I1 =>  inp_feat(263), I2 =>  inp_feat(306), I3 =>  inp_feat(375), I4 =>  inp_feat(215), I5 =>  inp_feat(186)); 
C_12_S_3_L_5_inst : LUT6 generic map(INIT => "0010001111000010100111110000101001001111111000000111111100000001") port map( O =>C_12_S_3_L_5_out, I0 =>  inp_feat(392), I1 =>  inp_feat(215), I2 =>  inp_feat(186), I3 =>  inp_feat(420), I4 =>  inp_feat(199), I5 =>  inp_feat(277)); 
C_12_S_4_L_0_inst : LUT6 generic map(INIT => "0001111110100101001001001010000110101010101000001011000011110010") port map( O =>C_12_S_4_L_0_out, I0 =>  inp_feat(372), I1 =>  inp_feat(233), I2 =>  inp_feat(374), I3 =>  inp_feat(417), I4 =>  inp_feat(149), I5 =>  inp_feat(485)); 
C_12_S_4_L_1_inst : LUT6 generic map(INIT => "1011000111101010111011000010000001001101000111101110111111000000") port map( O =>C_12_S_4_L_1_out, I0 =>  inp_feat(282), I1 =>  inp_feat(360), I2 =>  inp_feat(510), I3 =>  inp_feat(450), I4 =>  inp_feat(215), I5 =>  inp_feat(393)); 
C_12_S_4_L_2_inst : LUT6 generic map(INIT => "0000010100100000010010001101000011001001110000001100000011100100") port map( O =>C_12_S_4_L_2_out, I0 =>  inp_feat(250), I1 =>  inp_feat(289), I2 =>  inp_feat(296), I3 =>  inp_feat(186), I4 =>  inp_feat(215), I5 =>  inp_feat(393)); 
C_12_S_4_L_3_inst : LUT6 generic map(INIT => "1111101111011110101010110000101100000001000000001100111100000100") port map( O =>C_12_S_4_L_3_out, I0 =>  inp_feat(479), I1 =>  inp_feat(248), I2 =>  inp_feat(353), I3 =>  inp_feat(303), I4 =>  inp_feat(44), I5 =>  inp_feat(421)); 
C_12_S_4_L_4_inst : LUT6 generic map(INIT => "1010000001000100100100001111010100000000000011000010010001111100") port map( O =>C_12_S_4_L_4_out, I0 =>  inp_feat(17), I1 =>  inp_feat(452), I2 =>  inp_feat(375), I3 =>  inp_feat(496), I4 =>  inp_feat(440), I5 =>  inp_feat(490)); 
C_12_S_4_L_5_inst : LUT6 generic map(INIT => "0000011100000001011001110000011111111111000000110111111100010011") port map( O =>C_12_S_4_L_5_out, I0 =>  inp_feat(431), I1 =>  inp_feat(103), I2 =>  inp_feat(215), I3 =>  inp_feat(21), I4 =>  inp_feat(194), I5 =>  inp_feat(467)); 
C_12_S_5_L_0_inst : LUT6 generic map(INIT => "0100011101000111100001111111111111011101011101110111111111111111") port map( O =>C_12_S_5_L_0_out, I0 =>  inp_feat(126), I1 =>  inp_feat(306), I2 =>  inp_feat(417), I3 =>  inp_feat(186), I4 =>  inp_feat(215), I5 =>  inp_feat(103)); 
C_12_S_5_L_1_inst : LUT6 generic map(INIT => "0011010011100010101010100000000011100001100000001111111010100010") port map( O =>C_12_S_5_L_1_out, I0 =>  inp_feat(70), I1 =>  inp_feat(330), I2 =>  inp_feat(447), I3 =>  inp_feat(344), I4 =>  inp_feat(448), I5 =>  inp_feat(357)); 
C_12_S_5_L_2_inst : LUT6 generic map(INIT => "1101111000000010000101010000011111000101000000001110111000000000") port map( O =>C_12_S_5_L_2_out, I0 =>  inp_feat(368), I1 =>  inp_feat(308), I2 =>  inp_feat(446), I3 =>  inp_feat(402), I4 =>  inp_feat(215), I5 =>  inp_feat(211)); 
C_12_S_5_L_3_inst : LUT6 generic map(INIT => "0111100000110010001110000101000010101010000110001110111100001100") port map( O =>C_12_S_5_L_3_out, I0 =>  inp_feat(449), I1 =>  inp_feat(43), I2 =>  inp_feat(233), I3 =>  inp_feat(474), I4 =>  inp_feat(199), I5 =>  inp_feat(277)); 
C_12_S_5_L_4_inst : LUT6 generic map(INIT => "0011001000100010000000000001011111010000001001101100010101001111") port map( O =>C_12_S_5_L_4_out, I0 =>  inp_feat(222), I1 =>  inp_feat(353), I2 =>  inp_feat(226), I3 =>  inp_feat(117), I4 =>  inp_feat(444), I5 =>  inp_feat(140)); 
C_12_S_5_L_5_inst : LUT6 generic map(INIT => "1001100110111000010111101010100011111111110100101110001011101010") port map( O =>C_12_S_5_L_5_out, I0 =>  inp_feat(225), I1 =>  inp_feat(53), I2 =>  inp_feat(405), I3 =>  inp_feat(215), I4 =>  inp_feat(186), I5 =>  inp_feat(29)); 
C_13_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000001110001111100000101001111110111111111111111") port map( O =>C_13_S_0_L_0_out, I0 =>  inp_feat(194), I1 =>  inp_feat(306), I2 =>  inp_feat(392), I3 =>  inp_feat(108), I4 =>  inp_feat(248), I5 =>  inp_feat(239)); 
C_13_S_0_L_1_inst : LUT6 generic map(INIT => "1000010001010101000000010000000111111111111111110000000000000100") port map( O =>C_13_S_0_L_1_out, I0 =>  inp_feat(417), I1 =>  inp_feat(16), I2 =>  inp_feat(241), I3 =>  inp_feat(248), I4 =>  inp_feat(20), I5 =>  inp_feat(353)); 
C_13_S_0_L_2_inst : LUT6 generic map(INIT => "0000010100010010010001001111010100111000111100001111000111110001") port map( O =>C_13_S_0_L_2_out, I0 =>  inp_feat(392), I1 =>  inp_feat(472), I2 =>  inp_feat(206), I3 =>  inp_feat(149), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_13_S_0_L_3_inst : LUT6 generic map(INIT => "1110110101001000101111110000111100000000000000001001010100000000") port map( O =>C_13_S_0_L_3_out, I0 =>  inp_feat(38), I1 =>  inp_feat(356), I2 =>  inp_feat(180), I3 =>  inp_feat(0), I4 =>  inp_feat(429), I5 =>  inp_feat(428)); 
C_13_S_0_L_4_inst : LUT6 generic map(INIT => "0000110100000000000011000000010001101100000011001100111100001110") port map( O =>C_13_S_0_L_4_out, I0 =>  inp_feat(307), I1 =>  inp_feat(206), I2 =>  inp_feat(393), I3 =>  inp_feat(142), I4 =>  inp_feat(186), I5 =>  inp_feat(215)); 
C_13_S_0_L_5_inst : LUT6 generic map(INIT => "1110101010101100011011000000110000000100000010000000100010101000") port map( O =>C_13_S_0_L_5_out, I0 =>  inp_feat(208), I1 =>  inp_feat(65), I2 =>  inp_feat(215), I3 =>  inp_feat(235), I4 =>  inp_feat(113), I5 =>  inp_feat(285)); 
C_13_S_1_L_0_inst : LUT6 generic map(INIT => "1000010001010101000000010000000111111111111111110000000000000100") port map( O =>C_13_S_1_L_0_out, I0 =>  inp_feat(417), I1 =>  inp_feat(16), I2 =>  inp_feat(241), I3 =>  inp_feat(248), I4 =>  inp_feat(20), I5 =>  inp_feat(353)); 
C_13_S_1_L_1_inst : LUT6 generic map(INIT => "0000010100010010010001001111010100111000111100001111000111110001") port map( O =>C_13_S_1_L_1_out, I0 =>  inp_feat(392), I1 =>  inp_feat(472), I2 =>  inp_feat(206), I3 =>  inp_feat(149), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_13_S_1_L_2_inst : LUT6 generic map(INIT => "1110110101001000101111110000111100000000000000001001010100000000") port map( O =>C_13_S_1_L_2_out, I0 =>  inp_feat(38), I1 =>  inp_feat(356), I2 =>  inp_feat(180), I3 =>  inp_feat(0), I4 =>  inp_feat(429), I5 =>  inp_feat(428)); 
C_13_S_1_L_3_inst : LUT6 generic map(INIT => "0000110100000000000011000000010001101100000011001100111100001110") port map( O =>C_13_S_1_L_3_out, I0 =>  inp_feat(307), I1 =>  inp_feat(206), I2 =>  inp_feat(393), I3 =>  inp_feat(142), I4 =>  inp_feat(186), I5 =>  inp_feat(215)); 
C_13_S_1_L_4_inst : LUT6 generic map(INIT => "1110101010101100011011000000110000000100000010000000100010101000") port map( O =>C_13_S_1_L_4_out, I0 =>  inp_feat(208), I1 =>  inp_feat(65), I2 =>  inp_feat(215), I3 =>  inp_feat(235), I4 =>  inp_feat(113), I5 =>  inp_feat(285)); 
C_13_S_1_L_5_inst : LUT6 generic map(INIT => "0000000101010010001000000000100010000001100000111110110011100000") port map( O =>C_13_S_1_L_5_out, I0 =>  inp_feat(504), I1 =>  inp_feat(69), I2 =>  inp_feat(61), I3 =>  inp_feat(209), I4 =>  inp_feat(186), I5 =>  inp_feat(215)); 
C_13_S_2_L_0_inst : LUT6 generic map(INIT => "0000001011000100000011001111110100110110111001000100110011111111") port map( O =>C_13_S_2_L_0_out, I0 =>  inp_feat(393), I1 =>  inp_feat(257), I2 =>  inp_feat(476), I3 =>  inp_feat(199), I4 =>  inp_feat(353), I5 =>  inp_feat(334)); 
C_13_S_2_L_1_inst : LUT6 generic map(INIT => "1110100111010000000000001101000000100010000001000000000000000000") port map( O =>C_13_S_2_L_1_out, I0 =>  inp_feat(256), I1 =>  inp_feat(243), I2 =>  inp_feat(85), I3 =>  inp_feat(28), I4 =>  inp_feat(428), I5 =>  inp_feat(183)); 
C_13_S_2_L_2_inst : LUT6 generic map(INIT => "0001010100000111000000010100000011111111011111110000000100000010") port map( O =>C_13_S_2_L_2_out, I0 =>  inp_feat(149), I1 =>  inp_feat(403), I2 =>  inp_feat(123), I3 =>  inp_feat(429), I4 =>  inp_feat(428), I5 =>  inp_feat(417)); 
C_13_S_2_L_3_inst : LUT6 generic map(INIT => "1110011111110010100000101111000100100010111000010000000000001010") port map( O =>C_13_S_2_L_3_out, I0 =>  inp_feat(448), I1 =>  inp_feat(383), I2 =>  inp_feat(131), I3 =>  inp_feat(244), I4 =>  inp_feat(480), I5 =>  inp_feat(305)); 
C_13_S_2_L_4_inst : LUT6 generic map(INIT => "0001010100001000111010100000000001101000000010001111001100000000") port map( O =>C_13_S_2_L_4_out, I0 =>  inp_feat(250), I1 =>  inp_feat(239), I2 =>  inp_feat(24), I3 =>  inp_feat(301), I4 =>  inp_feat(186), I5 =>  inp_feat(215)); 
C_13_S_2_L_5_inst : LUT6 generic map(INIT => "1011111110100111100111110001011100000011000000110000010101100001") port map( O =>C_13_S_2_L_5_out, I0 =>  inp_feat(279), I1 =>  inp_feat(353), I2 =>  inp_feat(215), I3 =>  inp_feat(235), I4 =>  inp_feat(113), I5 =>  inp_feat(285)); 
C_13_S_3_L_0_inst : LUT6 generic map(INIT => "1000101011101100000010110100101100000000000100000000011001001011") port map( O =>C_13_S_3_L_0_out, I0 =>  inp_feat(117), I1 =>  inp_feat(128), I2 =>  inp_feat(176), I3 =>  inp_feat(353), I4 =>  inp_feat(31), I5 =>  inp_feat(301)); 
C_13_S_3_L_1_inst : LUT6 generic map(INIT => "0010100000001100101110000000000000000000000000000000000000000000") port map( O =>C_13_S_3_L_1_out, I0 =>  inp_feat(110), I1 =>  inp_feat(0), I2 =>  inp_feat(429), I3 =>  inp_feat(428), I4 =>  inp_feat(323), I5 =>  inp_feat(379)); 
C_13_S_3_L_2_inst : LUT6 generic map(INIT => "0000100011100000010011100000000010001100000000001100111100001100") port map( O =>C_13_S_3_L_2_out, I0 =>  inp_feat(494), I1 =>  inp_feat(276), I2 =>  inp_feat(241), I3 =>  inp_feat(484), I4 =>  inp_feat(121), I5 =>  inp_feat(122)); 
C_13_S_3_L_3_inst : LUT6 generic map(INIT => "0100111100011011000110010000010010100110100000000000000111000000") port map( O =>C_13_S_3_L_3_out, I0 =>  inp_feat(397), I1 =>  inp_feat(96), I2 =>  inp_feat(257), I3 =>  inp_feat(453), I4 =>  inp_feat(305), I5 =>  inp_feat(321)); 
C_13_S_3_L_4_inst : LUT6 generic map(INIT => "1111001100000011101001010000100000000000000100001000001010000000") port map( O =>C_13_S_3_L_4_out, I0 =>  inp_feat(413), I1 =>  inp_feat(239), I2 =>  inp_feat(369), I3 =>  inp_feat(152), I4 =>  inp_feat(21), I5 =>  inp_feat(221)); 
C_13_S_3_L_5_inst : LUT6 generic map(INIT => "0100010001000100010011001000110011011100000000001100111000000000") port map( O =>C_13_S_3_L_5_out, I0 =>  inp_feat(37), I1 =>  inp_feat(428), I2 =>  inp_feat(417), I3 =>  inp_feat(468), I4 =>  inp_feat(403), I5 =>  inp_feat(103)); 
C_13_S_4_L_0_inst : LUT6 generic map(INIT => "0101100100000011010100000000100110110011000000001111011000100000") port map( O =>C_13_S_4_L_0_out, I0 =>  inp_feat(440), I1 =>  inp_feat(279), I2 =>  inp_feat(349), I3 =>  inp_feat(428), I4 =>  inp_feat(149), I5 =>  inp_feat(211)); 
C_13_S_4_L_1_inst : LUT6 generic map(INIT => "1111101010011101000000000000110000000010100000010000000000000000") port map( O =>C_13_S_4_L_1_out, I0 =>  inp_feat(403), I1 =>  inp_feat(334), I2 =>  inp_feat(362), I3 =>  inp_feat(427), I4 =>  inp_feat(428), I5 =>  inp_feat(421)); 
C_13_S_4_L_2_inst : LUT6 generic map(INIT => "0001000100000011001000110111111111010111000111110011111111111111") port map( O =>C_13_S_4_L_2_out, I0 =>  inp_feat(180), I1 =>  inp_feat(123), I2 =>  inp_feat(353), I3 =>  inp_feat(199), I4 =>  inp_feat(417), I5 =>  inp_feat(277)); 
C_13_S_4_L_3_inst : LUT6 generic map(INIT => "1000011011000000000101100000001000001000000000001110000100000001") port map( O =>C_13_S_4_L_3_out, I0 =>  inp_feat(460), I1 =>  inp_feat(78), I2 =>  inp_feat(499), I3 =>  inp_feat(171), I4 =>  inp_feat(92), I5 =>  inp_feat(494)); 
C_13_S_4_L_4_inst : LUT6 generic map(INIT => "1011011100011111001101010001111101010111010011110110011111011101") port map( O =>C_13_S_4_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(190), I2 =>  inp_feat(403), I3 =>  inp_feat(103), I4 =>  inp_feat(233), I5 =>  inp_feat(263)); 
C_13_S_4_L_5_inst : LUT6 generic map(INIT => "0100010001010001010101000000100010010000000111001101100000000000") port map( O =>C_13_S_4_L_5_out, I0 =>  inp_feat(244), I1 =>  inp_feat(509), I2 =>  inp_feat(43), I3 =>  inp_feat(483), I4 =>  inp_feat(152), I5 =>  inp_feat(358)); 
C_13_S_5_L_0_inst : LUT6 generic map(INIT => "0110111010100100010101001000110011001100000011000000110000001000") port map( O =>C_13_S_5_L_0_out, I0 =>  inp_feat(417), I1 =>  inp_feat(225), I2 =>  inp_feat(126), I3 =>  inp_feat(95), I4 =>  inp_feat(439), I5 =>  inp_feat(323)); 
C_13_S_5_L_1_inst : LUT6 generic map(INIT => "1011000010010011111111100000110000001000011110010000000010000000") port map( O =>C_13_S_5_L_1_out, I0 =>  inp_feat(446), I1 =>  inp_feat(404), I2 =>  inp_feat(25), I3 =>  inp_feat(299), I4 =>  inp_feat(263), I5 =>  inp_feat(305)); 
C_13_S_5_L_2_inst : LUT6 generic map(INIT => "0101001000010001110011010110000000000010000000000100100001100000") port map( O =>C_13_S_5_L_2_out, I0 =>  inp_feat(108), I1 =>  inp_feat(92), I2 =>  inp_feat(404), I3 =>  inp_feat(484), I4 =>  inp_feat(229), I5 =>  inp_feat(494)); 
C_13_S_5_L_3_inst : LUT6 generic map(INIT => "1101010010000000010111000000000000011100000000000000000000001000") port map( O =>C_13_S_5_L_3_out, I0 =>  inp_feat(322), I1 =>  inp_feat(196), I2 =>  inp_feat(330), I3 =>  inp_feat(56), I4 =>  inp_feat(171), I5 =>  inp_feat(494)); 
C_13_S_5_L_4_inst : LUT6 generic map(INIT => "0110001011110000000001101100010000000100110000100000000000000000") port map( O =>C_13_S_5_L_4_out, I0 =>  inp_feat(362), I1 =>  inp_feat(194), I2 =>  inp_feat(193), I3 =>  inp_feat(175), I4 =>  inp_feat(428), I5 =>  inp_feat(421)); 
C_13_S_5_L_5_inst : LUT6 generic map(INIT => "1100001110010001110101110001011100010001000010010101000100010101") port map( O =>C_13_S_5_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(248), I2 =>  inp_feat(282), I3 =>  inp_feat(71), I4 =>  inp_feat(510), I5 =>  inp_feat(220)); 
C_14_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000110001111100000100001111110101111111111111") port map( O =>C_14_S_0_L_0_out, I0 =>  inp_feat(353), I1 =>  inp_feat(306), I2 =>  inp_feat(392), I3 =>  inp_feat(108), I4 =>  inp_feat(248), I5 =>  inp_feat(239)); 
C_14_S_0_L_1_inst : LUT6 generic map(INIT => "0000110000000110101000100000001000101111000000111011111010100000") port map( O =>C_14_S_0_L_1_out, I0 =>  inp_feat(386), I1 =>  inp_feat(190), I2 =>  inp_feat(82), I3 =>  inp_feat(51), I4 =>  inp_feat(215), I5 =>  inp_feat(431)); 
C_14_S_0_L_2_inst : LUT6 generic map(INIT => "1110111011100000111011100110001011000000111000101011001011111011") port map( O =>C_14_S_0_L_2_out, I0 =>  inp_feat(257), I1 =>  inp_feat(248), I2 =>  inp_feat(48), I3 =>  inp_feat(352), I4 =>  inp_feat(199), I5 =>  inp_feat(353)); 
C_14_S_0_L_3_inst : LUT6 generic map(INIT => "0000000100000111111001111101111110101010101101111011111111111111") port map( O =>C_14_S_0_L_3_out, I0 =>  inp_feat(239), I1 =>  inp_feat(393), I2 =>  inp_feat(279), I3 =>  inp_feat(352), I4 =>  inp_feat(199), I5 =>  inp_feat(353)); 
C_14_S_0_L_4_inst : LUT6 generic map(INIT => "1001000000000000011111010010000011010110000000001111111110000000") port map( O =>C_14_S_0_L_4_out, I0 =>  inp_feat(215), I1 =>  inp_feat(431), I2 =>  inp_feat(345), I3 =>  inp_feat(314), I4 =>  inp_feat(186), I5 =>  inp_feat(194)); 
C_14_S_0_L_5_inst : LUT6 generic map(INIT => "1010000000000001101100100000001000000000000000000111000000000010") port map( O =>C_14_S_0_L_5_out, I0 =>  inp_feat(145), I1 =>  inp_feat(509), I2 =>  inp_feat(64), I3 =>  inp_feat(366), I4 =>  inp_feat(61), I5 =>  inp_feat(85)); 
C_14_S_1_L_0_inst : LUT6 generic map(INIT => "0000110000000110101000100000001000101111000000111011111010100000") port map( O =>C_14_S_1_L_0_out, I0 =>  inp_feat(386), I1 =>  inp_feat(190), I2 =>  inp_feat(82), I3 =>  inp_feat(51), I4 =>  inp_feat(215), I5 =>  inp_feat(431)); 
C_14_S_1_L_1_inst : LUT6 generic map(INIT => "1110111011100000111011100110001011000000111000101011001011111011") port map( O =>C_14_S_1_L_1_out, I0 =>  inp_feat(257), I1 =>  inp_feat(248), I2 =>  inp_feat(48), I3 =>  inp_feat(352), I4 =>  inp_feat(199), I5 =>  inp_feat(353)); 
C_14_S_1_L_2_inst : LUT6 generic map(INIT => "0000000100000111111001111101111110101010101101111011111111111111") port map( O =>C_14_S_1_L_2_out, I0 =>  inp_feat(239), I1 =>  inp_feat(393), I2 =>  inp_feat(279), I3 =>  inp_feat(352), I4 =>  inp_feat(199), I5 =>  inp_feat(353)); 
C_14_S_1_L_3_inst : LUT6 generic map(INIT => "1001000000000000011111010010000011010110000000001111111110000000") port map( O =>C_14_S_1_L_3_out, I0 =>  inp_feat(215), I1 =>  inp_feat(431), I2 =>  inp_feat(345), I3 =>  inp_feat(314), I4 =>  inp_feat(186), I5 =>  inp_feat(194)); 
C_14_S_1_L_4_inst : LUT6 generic map(INIT => "1010000000000001101100100000001000000000000000000111000000000010") port map( O =>C_14_S_1_L_4_out, I0 =>  inp_feat(145), I1 =>  inp_feat(509), I2 =>  inp_feat(64), I3 =>  inp_feat(366), I4 =>  inp_feat(61), I5 =>  inp_feat(85)); 
C_14_S_1_L_5_inst : LUT6 generic map(INIT => "0001110100000000010111000000001011001100000100001101111100000100") port map( O =>C_14_S_1_L_5_out, I0 =>  inp_feat(431), I1 =>  inp_feat(363), I2 =>  inp_feat(461), I3 =>  inp_feat(76), I4 =>  inp_feat(194), I5 =>  inp_feat(485)); 
C_14_S_2_L_0_inst : LUT6 generic map(INIT => "1101000001110101011100111111111111110001111101111111011111111111") port map( O =>C_14_S_2_L_0_out, I0 =>  inp_feat(431), I1 =>  inp_feat(103), I2 =>  inp_feat(391), I3 =>  inp_feat(215), I4 =>  inp_feat(393), I5 =>  inp_feat(497)); 
C_14_S_2_L_1_inst : LUT6 generic map(INIT => "0000000000001010101000101110100010010000110001001000100011101010") port map( O =>C_14_S_2_L_1_out, I0 =>  inp_feat(460), I1 =>  inp_feat(379), I2 =>  inp_feat(363), I3 =>  inp_feat(417), I4 =>  inp_feat(194), I5 =>  inp_feat(485)); 
C_14_S_2_L_2_inst : LUT6 generic map(INIT => "0010101100011110011100111011110000000000000010001010111000000000") port map( O =>C_14_S_2_L_2_out, I0 =>  inp_feat(210), I1 =>  inp_feat(115), I2 =>  inp_feat(445), I3 =>  inp_feat(389), I4 =>  inp_feat(61), I5 =>  inp_feat(85)); 
C_14_S_2_L_3_inst : LUT6 generic map(INIT => "1111001011111110111100110011000100010000000000100000000001110000") port map( O =>C_14_S_2_L_3_out, I0 =>  inp_feat(510), I1 =>  inp_feat(47), I2 =>  inp_feat(384), I3 =>  inp_feat(27), I4 =>  inp_feat(394), I5 =>  inp_feat(370)); 
C_14_S_2_L_4_inst : LUT6 generic map(INIT => "1100000100001000010010000000000000000001000000000000000000000100") port map( O =>C_14_S_2_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(375), I2 =>  inp_feat(355), I3 =>  inp_feat(77), I4 =>  inp_feat(387), I5 =>  inp_feat(76)); 
C_14_S_2_L_5_inst : LUT6 generic map(INIT => "0101001001100010010100100000001000000000000000000000000001000000") port map( O =>C_14_S_2_L_5_out, I0 =>  inp_feat(186), I1 =>  inp_feat(409), I2 =>  inp_feat(291), I3 =>  inp_feat(119), I4 =>  inp_feat(109), I5 =>  inp_feat(314)); 
C_14_S_3_L_0_inst : LUT6 generic map(INIT => "1101100001110101010100011111111111000001111101111111011111111111") port map( O =>C_14_S_3_L_0_out, I0 =>  inp_feat(431), I1 =>  inp_feat(103), I2 =>  inp_feat(391), I3 =>  inp_feat(215), I4 =>  inp_feat(393), I5 =>  inp_feat(497)); 
C_14_S_3_L_1_inst : LUT6 generic map(INIT => "0001111000010000000110001111010001011000011100011111000011110011") port map( O =>C_14_S_3_L_1_out, I0 =>  inp_feat(126), I1 =>  inp_feat(199), I2 =>  inp_feat(350), I3 =>  inp_feat(393), I4 =>  inp_feat(215), I5 =>  inp_feat(103)); 
C_14_S_3_L_2_inst : LUT6 generic map(INIT => "0001000011000000100111010000000011111110100000001100110101001100") port map( O =>C_14_S_3_L_2_out, I0 =>  inp_feat(75), I1 =>  inp_feat(371), I2 =>  inp_feat(227), I3 =>  inp_feat(237), I4 =>  inp_feat(186), I5 =>  inp_feat(403)); 
C_14_S_3_L_3_inst : LUT6 generic map(INIT => "1000010011000101000101000000010000000000000000000000000001000001") port map( O =>C_14_S_3_L_3_out, I0 =>  inp_feat(211), I1 =>  inp_feat(432), I2 =>  inp_feat(194), I3 =>  inp_feat(235), I4 =>  inp_feat(109), I5 =>  inp_feat(314)); 
C_14_S_3_L_4_inst : LUT6 generic map(INIT => "1101110100010001011000101101011000000001000000000011000100001000") port map( O =>C_14_S_3_L_4_out, I0 =>  inp_feat(39), I1 =>  inp_feat(221), I2 =>  inp_feat(454), I3 =>  inp_feat(449), I4 =>  inp_feat(299), I5 =>  inp_feat(85)); 
C_14_S_3_L_5_inst : LUT6 generic map(INIT => "0100000010001101011011110000100000000000000001001000110000000000") port map( O =>C_14_S_3_L_5_out, I0 =>  inp_feat(181), I1 =>  inp_feat(366), I2 =>  inp_feat(306), I3 =>  inp_feat(265), I4 =>  inp_feat(299), I5 =>  inp_feat(85)); 
C_14_S_4_L_0_inst : LUT6 generic map(INIT => "1110100100001100000000001110010000000000000010000000000011010000") port map( O =>C_14_S_4_L_0_out, I0 =>  inp_feat(208), I1 =>  inp_feat(370), I2 =>  inp_feat(235), I3 =>  inp_feat(468), I4 =>  inp_feat(372), I5 =>  inp_feat(237)); 
C_14_S_4_L_1_inst : LUT6 generic map(INIT => "0000110111010100000001000001010011011111000000010000000000000100") port map( O =>C_14_S_4_L_1_out, I0 =>  inp_feat(367), I1 =>  inp_feat(224), I2 =>  inp_feat(267), I3 =>  inp_feat(506), I4 =>  inp_feat(507), I5 =>  inp_feat(400)); 
C_14_S_4_L_2_inst : LUT6 generic map(INIT => "0000110110010011110000011000000000000101110110111110100010000000") port map( O =>C_14_S_4_L_2_out, I0 =>  inp_feat(350), I1 =>  inp_feat(115), I2 =>  inp_feat(61), I3 =>  inp_feat(376), I4 =>  inp_feat(215), I5 =>  inp_feat(121)); 
C_14_S_4_L_3_inst : LUT6 generic map(INIT => "1111101010100001000000001110000000010001000000100000000000000000") port map( O =>C_14_S_4_L_3_out, I0 =>  inp_feat(387), I1 =>  inp_feat(110), I2 =>  inp_feat(232), I3 =>  inp_feat(5), I4 =>  inp_feat(67), I5 =>  inp_feat(366)); 
C_14_S_4_L_4_inst : LUT6 generic map(INIT => "0111000010010000000011000000100000001101001110001010110001111000") port map( O =>C_14_S_4_L_4_out, I0 =>  inp_feat(175), I1 =>  inp_feat(222), I2 =>  inp_feat(279), I3 =>  inp_feat(294), I4 =>  inp_feat(497), I5 =>  inp_feat(121)); 
C_14_S_4_L_5_inst : LUT6 generic map(INIT => "0111000110000001100100010100000011111111001110000001000100000001") port map( O =>C_14_S_4_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(393), I2 =>  inp_feat(43), I3 =>  inp_feat(376), I4 =>  inp_feat(139), I5 =>  inp_feat(306)); 
C_14_S_5_L_0_inst : LUT6 generic map(INIT => "0000001010101011000000100010001110001011000101110000000000100000") port map( O =>C_14_S_5_L_0_out, I0 =>  inp_feat(296), I1 =>  inp_feat(254), I2 =>  inp_feat(48), I3 =>  inp_feat(12), I4 =>  inp_feat(507), I5 =>  inp_feat(400)); 
C_14_S_5_L_1_inst : LUT6 generic map(INIT => "1000001110011111001101111111111110111101000010110111111111111111") port map( O =>C_14_S_5_L_1_out, I0 =>  inp_feat(353), I1 =>  inp_feat(215), I2 =>  inp_feat(306), I3 =>  inp_feat(321), I4 =>  inp_feat(393), I5 =>  inp_feat(497)); 
C_14_S_5_L_2_inst : LUT6 generic map(INIT => "0000001100001000010000001100110011000000100100001100000011001100") port map( O =>C_14_S_5_L_2_out, I0 =>  inp_feat(413), I1 =>  inp_feat(165), I2 =>  inp_feat(14), I3 =>  inp_feat(353), I4 =>  inp_feat(352), I5 =>  inp_feat(306)); 
C_14_S_5_L_3_inst : LUT6 generic map(INIT => "0010000010100010101110011011010111010010011000001011000000000000") port map( O =>C_14_S_5_L_3_out, I0 =>  inp_feat(206), I1 =>  inp_feat(47), I2 =>  inp_feat(162), I3 =>  inp_feat(438), I4 =>  inp_feat(467), I5 =>  inp_feat(405)); 
C_14_S_5_L_4_inst : LUT6 generic map(INIT => "1101110101110111100000011011001100010101001100011101000100010001") port map( O =>C_14_S_5_L_4_out, I0 =>  inp_feat(215), I1 =>  inp_feat(186), I2 =>  inp_feat(92), I3 =>  inp_feat(194), I4 =>  inp_feat(261), I5 =>  inp_feat(482)); 
C_14_S_5_L_5_inst : LUT6 generic map(INIT => "0000010001000000000100010011000010011100000011000000000000000000") port map( O =>C_14_S_5_L_5_out, I0 =>  inp_feat(37), I1 =>  inp_feat(158), I2 =>  inp_feat(327), I3 =>  inp_feat(466), I4 =>  inp_feat(2), I5 =>  inp_feat(8)); 
C_15_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000100110101111100000100011111110111111111111111") port map( O =>C_15_S_0_L_0_out, I0 =>  inp_feat(279), I1 =>  inp_feat(306), I2 =>  inp_feat(392), I3 =>  inp_feat(108), I4 =>  inp_feat(248), I5 =>  inp_feat(239)); 
C_15_S_0_L_1_inst : LUT6 generic map(INIT => "0101010100000000111111110001000011110111000000001111111100001001") port map( O =>C_15_S_0_L_1_out, I0 =>  inp_feat(199), I1 =>  inp_feat(180), I2 =>  inp_feat(395), I3 =>  inp_feat(312), I4 =>  inp_feat(186), I5 =>  inp_feat(445)); 
C_15_S_0_L_2_inst : LUT6 generic map(INIT => "1110001001000100111110000000100010101100000011001100100010000000") port map( O =>C_15_S_0_L_2_out, I0 =>  inp_feat(142), I1 =>  inp_feat(225), I2 =>  inp_feat(224), I3 =>  inp_feat(98), I4 =>  inp_feat(239), I5 =>  inp_feat(7)); 
C_15_S_0_L_3_inst : LUT6 generic map(INIT => "0001000010000001110111100000100010111010000000101000101000001000") port map( O =>C_15_S_0_L_3_out, I0 =>  inp_feat(115), I1 =>  inp_feat(460), I2 =>  inp_feat(445), I3 =>  inp_feat(28), I4 =>  inp_feat(239), I5 =>  inp_feat(7)); 
C_15_S_0_L_4_inst : LUT6 generic map(INIT => "0010110001100110010001011101110111001100010011101110111011011111") port map( O =>C_15_S_0_L_4_out, I0 =>  inp_feat(190), I1 =>  inp_feat(387), I2 =>  inp_feat(173), I3 =>  inp_feat(403), I4 =>  inp_feat(186), I5 =>  inp_feat(485)); 
C_15_S_0_L_5_inst : LUT6 generic map(INIT => "0100010011001101101110000100110000101100110011001011001001000110") port map( O =>C_15_S_0_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(50), I2 =>  inp_feat(417), I3 =>  inp_feat(393), I4 =>  inp_feat(224), I5 =>  inp_feat(440)); 
C_15_S_1_L_0_inst : LUT6 generic map(INIT => "0101010100000000111111110001000011110111000000001111111100001001") port map( O =>C_15_S_1_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(180), I2 =>  inp_feat(395), I3 =>  inp_feat(312), I4 =>  inp_feat(186), I5 =>  inp_feat(445)); 
C_15_S_1_L_1_inst : LUT6 generic map(INIT => "1110001001000100111110000000100010101100000011001100100010000000") port map( O =>C_15_S_1_L_1_out, I0 =>  inp_feat(142), I1 =>  inp_feat(225), I2 =>  inp_feat(224), I3 =>  inp_feat(98), I4 =>  inp_feat(239), I5 =>  inp_feat(7)); 
C_15_S_1_L_2_inst : LUT6 generic map(INIT => "0001000010000001110111100000100010111010000000101000101000001000") port map( O =>C_15_S_1_L_2_out, I0 =>  inp_feat(115), I1 =>  inp_feat(460), I2 =>  inp_feat(445), I3 =>  inp_feat(28), I4 =>  inp_feat(239), I5 =>  inp_feat(7)); 
C_15_S_1_L_3_inst : LUT6 generic map(INIT => "0010110001100110010001011101110111001100010011101110111011011111") port map( O =>C_15_S_1_L_3_out, I0 =>  inp_feat(190), I1 =>  inp_feat(387), I2 =>  inp_feat(173), I3 =>  inp_feat(403), I4 =>  inp_feat(186), I5 =>  inp_feat(485)); 
C_15_S_1_L_4_inst : LUT6 generic map(INIT => "0100010011001101101110000100110000101100110011001011001001000110") port map( O =>C_15_S_1_L_4_out, I0 =>  inp_feat(215), I1 =>  inp_feat(50), I2 =>  inp_feat(417), I3 =>  inp_feat(393), I4 =>  inp_feat(224), I5 =>  inp_feat(440)); 
C_15_S_1_L_5_inst : LUT6 generic map(INIT => "1011111011010100110111000000000010111011000111110000000000000000") port map( O =>C_15_S_1_L_5_out, I0 =>  inp_feat(84), I1 =>  inp_feat(368), I2 =>  inp_feat(445), I3 =>  inp_feat(216), I4 =>  inp_feat(94), I5 =>  inp_feat(381)); 
C_15_S_2_L_0_inst : LUT6 generic map(INIT => "0100101000001000110010000001100010001100000010001010101000001000") port map( O =>C_15_S_2_L_0_out, I0 =>  inp_feat(207), I1 =>  inp_feat(98), I2 =>  inp_feat(445), I3 =>  inp_feat(28), I4 =>  inp_feat(194), I5 =>  inp_feat(239)); 
C_15_S_2_L_1_inst : LUT6 generic map(INIT => "1001010100000000011110110011000011111011000100001111111101110000") port map( O =>C_15_S_2_L_1_out, I0 =>  inp_feat(190), I1 =>  inp_feat(239), I2 =>  inp_feat(24), I3 =>  inp_feat(28), I4 =>  inp_feat(215), I5 =>  inp_feat(211)); 
C_15_S_2_L_2_inst : LUT6 generic map(INIT => "0011000100011001101000000000000011111001001110011010100000001000") port map( O =>C_15_S_2_L_2_out, I0 =>  inp_feat(96), I1 =>  inp_feat(316), I2 =>  inp_feat(436), I3 =>  inp_feat(453), I4 =>  inp_feat(186), I5 =>  inp_feat(215)); 
C_15_S_2_L_3_inst : LUT6 generic map(INIT => "1101110111101101101010101000000011101101111000011000100011000000") port map( O =>C_15_S_2_L_3_out, I0 =>  inp_feat(344), I1 =>  inp_feat(77), I2 =>  inp_feat(404), I3 =>  inp_feat(313), I4 =>  inp_feat(181), I5 =>  inp_feat(440)); 
C_15_S_2_L_4_inst : LUT6 generic map(INIT => "0000010000010101111110001001000011011111000011111111000000000000") port map( O =>C_15_S_2_L_4_out, I0 =>  inp_feat(476), I1 =>  inp_feat(332), I2 =>  inp_feat(17), I3 =>  inp_feat(361), I4 =>  inp_feat(485), I5 =>  inp_feat(440)); 
C_15_S_2_L_5_inst : LUT6 generic map(INIT => "1011111000011101100100000000110010000000000001000000000000000000") port map( O =>C_15_S_2_L_5_out, I0 =>  inp_feat(239), I1 =>  inp_feat(361), I2 =>  inp_feat(353), I3 =>  inp_feat(445), I4 =>  inp_feat(197), I5 =>  inp_feat(145)); 
C_15_S_3_L_0_inst : LUT6 generic map(INIT => "0100100100001100001111001000110010111000111010001100111011001100") port map( O =>C_15_S_3_L_0_out, I0 =>  inp_feat(483), I1 =>  inp_feat(46), I2 =>  inp_feat(91), I3 =>  inp_feat(215), I4 =>  inp_feat(211), I5 =>  inp_feat(489)); 
C_15_S_3_L_1_inst : LUT6 generic map(INIT => "1000101000101000101101010101000111011001001000101111011101110000") port map( O =>C_15_S_3_L_1_out, I0 =>  inp_feat(239), I1 =>  inp_feat(103), I2 =>  inp_feat(24), I3 =>  inp_feat(28), I4 =>  inp_feat(215), I5 =>  inp_feat(431)); 
C_15_S_3_L_2_inst : LUT6 generic map(INIT => "0100000010100000110111010101000111111001001000101111011101110000") port map( O =>C_15_S_3_L_2_out, I0 =>  inp_feat(239), I1 =>  inp_feat(103), I2 =>  inp_feat(24), I3 =>  inp_feat(28), I4 =>  inp_feat(215), I5 =>  inp_feat(431)); 
C_15_S_3_L_3_inst : LUT6 generic map(INIT => "1101011111111111000000110000100011010011001100111000110010000100") port map( O =>C_15_S_3_L_3_out, I0 =>  inp_feat(123), I1 =>  inp_feat(239), I2 =>  inp_feat(199), I3 =>  inp_feat(344), I4 =>  inp_feat(50), I5 =>  inp_feat(176)); 
C_15_S_3_L_4_inst : LUT6 generic map(INIT => "0001100001111111000100110111111111101000011001110001011111111111") port map( O =>C_15_S_3_L_4_out, I0 =>  inp_feat(186), I1 =>  inp_feat(334), I2 =>  inp_feat(123), I3 =>  inp_feat(215), I4 =>  inp_feat(510), I5 =>  inp_feat(7)); 
C_15_S_3_L_5_inst : LUT6 generic map(INIT => "1111101011110101000100011101000111111100001111010000000000000000") port map( O =>C_15_S_3_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(239), I2 =>  inp_feat(21), I3 =>  inp_feat(467), I4 =>  inp_feat(94), I5 =>  inp_feat(381)); 
C_15_S_4_L_0_inst : LUT6 generic map(INIT => "1010100000011000101010000000100011011100100010001111111011100010") port map( O =>C_15_S_4_L_0_out, I0 =>  inp_feat(168), I1 =>  inp_feat(378), I2 =>  inp_feat(262), I3 =>  inp_feat(28), I4 =>  inp_feat(194), I5 =>  inp_feat(239)); 
C_15_S_4_L_1_inst : LUT6 generic map(INIT => "0100000110111000000000000010000010101100101010000000100011000010") port map( O =>C_15_S_4_L_1_out, I0 =>  inp_feat(142), I1 =>  inp_feat(136), I2 =>  inp_feat(510), I3 =>  inp_feat(370), I4 =>  inp_feat(285), I5 =>  inp_feat(467)); 
C_15_S_4_L_2_inst : LUT6 generic map(INIT => "1010101011000010100010111000001100100001010010000000000001000000") port map( O =>C_15_S_4_L_2_out, I0 =>  inp_feat(140), I1 =>  inp_feat(395), I2 =>  inp_feat(179), I3 =>  inp_feat(309), I4 =>  inp_feat(419), I5 =>  inp_feat(312)); 
C_15_S_4_L_3_inst : LUT6 generic map(INIT => "0001000100000001110110000000000011111001000010100000000000000000") port map( O =>C_15_S_4_L_3_out, I0 =>  inp_feat(269), I1 =>  inp_feat(368), I2 =>  inp_feat(445), I3 =>  inp_feat(216), I4 =>  inp_feat(94), I5 =>  inp_feat(381)); 
C_15_S_4_L_4_inst : LUT6 generic map(INIT => "1101101111101000001111000001001000010001101110000000000000000000") port map( O =>C_15_S_4_L_4_out, I0 =>  inp_feat(368), I1 =>  inp_feat(291), I2 =>  inp_feat(379), I3 =>  inp_feat(243), I4 =>  inp_feat(398), I5 =>  inp_feat(107)); 
C_15_S_4_L_5_inst : LUT6 generic map(INIT => "0101010000000111100001010000000010000100110000001111001000000000") port map( O =>C_15_S_4_L_5_out, I0 =>  inp_feat(248), I1 =>  inp_feat(308), I2 =>  inp_feat(355), I3 =>  inp_feat(4), I4 =>  inp_feat(329), I5 =>  inp_feat(276)); 
C_15_S_5_L_0_inst : LUT6 generic map(INIT => "1010001100111111000101111101111101000001010011110000001000100001") port map( O =>C_15_S_5_L_0_out, I0 =>  inp_feat(392), I1 =>  inp_feat(170), I2 =>  inp_feat(215), I3 =>  inp_feat(211), I4 =>  inp_feat(480), I5 =>  inp_feat(265)); 
C_15_S_5_L_1_inst : LUT6 generic map(INIT => "1101111101011111000100100011000000000101000111010000101010100010") port map( O =>C_15_S_5_L_1_out, I0 =>  inp_feat(353), I1 =>  inp_feat(243), I2 =>  inp_feat(182), I3 =>  inp_feat(29), I4 =>  inp_feat(191), I5 =>  inp_feat(100)); 
C_15_S_5_L_2_inst : LUT6 generic map(INIT => "1000000010101100000000001010010100000010101000100000000000000000") port map( O =>C_15_S_5_L_2_out, I0 =>  inp_feat(228), I1 =>  inp_feat(475), I2 =>  inp_feat(191), I3 =>  inp_feat(288), I4 =>  inp_feat(274), I5 =>  inp_feat(378)); 
C_15_S_5_L_3_inst : LUT6 generic map(INIT => "0001000100000000000100010000010011110011000100000001000100000000") port map( O =>C_15_S_5_L_3_out, I0 =>  inp_feat(186), I1 =>  inp_feat(445), I2 =>  inp_feat(461), I3 =>  inp_feat(212), I4 =>  inp_feat(112), I5 =>  inp_feat(29)); 
C_15_S_5_L_4_inst : LUT6 generic map(INIT => "1101010111010110111000110011000001101010110000010000000000000000") port map( O =>C_15_S_5_L_4_out, I0 =>  inp_feat(415), I1 =>  inp_feat(322), I2 =>  inp_feat(407), I3 =>  inp_feat(111), I4 =>  inp_feat(128), I5 =>  inp_feat(400)); 
C_15_S_5_L_5_inst : LUT6 generic map(INIT => "0110111000100000000010011011011011110100000010000011101010110010") port map( O =>C_15_S_5_L_5_out, I0 =>  inp_feat(160), I1 =>  inp_feat(205), I2 =>  inp_feat(289), I3 =>  inp_feat(164), I4 =>  inp_feat(130), I5 =>  inp_feat(313)); 
C_16_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000110001111100000100001111110101111111111111") port map( O =>C_16_S_0_L_0_out, I0 =>  inp_feat(353), I1 =>  inp_feat(306), I2 =>  inp_feat(392), I3 =>  inp_feat(108), I4 =>  inp_feat(248), I5 =>  inp_feat(239)); 
C_16_S_0_L_1_inst : LUT6 generic map(INIT => "0001000110110001011110010001000001110011101100011111010101110000") port map( O =>C_16_S_0_L_1_out, I0 =>  inp_feat(393), I1 =>  inp_feat(215), I2 =>  inp_feat(78), I3 =>  inp_feat(210), I4 =>  inp_feat(227), I5 =>  inp_feat(497)); 
C_16_S_0_L_2_inst : LUT6 generic map(INIT => "1000011100000000100000101100000010001000110110001100000011101000") port map( O =>C_16_S_0_L_2_out, I0 =>  inp_feat(304), I1 =>  inp_feat(312), I2 =>  inp_feat(420), I3 =>  inp_feat(445), I4 =>  inp_feat(279), I5 =>  inp_feat(263)); 
C_16_S_0_L_3_inst : LUT6 generic map(INIT => "0010011000001100010111001100110001101110010111010111110111011101") port map( O =>C_16_S_0_L_3_out, I0 =>  inp_feat(194), I1 =>  inp_feat(214), I2 =>  inp_feat(199), I3 =>  inp_feat(403), I4 =>  inp_feat(103), I5 =>  inp_feat(485)); 
C_16_S_0_L_4_inst : LUT6 generic map(INIT => "0001111100001000101101110001101011110111000110000111010100000000") port map( O =>C_16_S_0_L_4_out, I0 =>  inp_feat(215), I1 =>  inp_feat(186), I2 =>  inp_feat(487), I3 =>  inp_feat(20), I4 =>  inp_feat(339), I5 =>  inp_feat(510)); 
C_16_S_0_L_5_inst : LUT6 generic map(INIT => "1100010111111000100000001010000011110001001110101000000010101100") port map( O =>C_16_S_0_L_5_out, I0 =>  inp_feat(386), I1 =>  inp_feat(452), I2 =>  inp_feat(20), I3 =>  inp_feat(445), I4 =>  inp_feat(393), I5 =>  inp_feat(456)); 
C_16_S_1_L_0_inst : LUT6 generic map(INIT => "0001000110110001011110010001000001110011101100011111010101110000") port map( O =>C_16_S_1_L_0_out, I0 =>  inp_feat(393), I1 =>  inp_feat(215), I2 =>  inp_feat(78), I3 =>  inp_feat(210), I4 =>  inp_feat(227), I5 =>  inp_feat(497)); 
C_16_S_1_L_1_inst : LUT6 generic map(INIT => "1000011100000000100000101100000010001000110110001100000011101000") port map( O =>C_16_S_1_L_1_out, I0 =>  inp_feat(304), I1 =>  inp_feat(312), I2 =>  inp_feat(420), I3 =>  inp_feat(445), I4 =>  inp_feat(279), I5 =>  inp_feat(263)); 
C_16_S_1_L_2_inst : LUT6 generic map(INIT => "0010011000001100010111001100110001101110010111010111110111011101") port map( O =>C_16_S_1_L_2_out, I0 =>  inp_feat(194), I1 =>  inp_feat(214), I2 =>  inp_feat(199), I3 =>  inp_feat(403), I4 =>  inp_feat(103), I5 =>  inp_feat(485)); 
C_16_S_1_L_3_inst : LUT6 generic map(INIT => "0001111100001000101101110001101011110111000110000111010100000000") port map( O =>C_16_S_1_L_3_out, I0 =>  inp_feat(215), I1 =>  inp_feat(186), I2 =>  inp_feat(487), I3 =>  inp_feat(20), I4 =>  inp_feat(339), I5 =>  inp_feat(510)); 
C_16_S_1_L_4_inst : LUT6 generic map(INIT => "1100010111111000100000001010000011110001001110101000000010101100") port map( O =>C_16_S_1_L_4_out, I0 =>  inp_feat(386), I1 =>  inp_feat(452), I2 =>  inp_feat(20), I3 =>  inp_feat(445), I4 =>  inp_feat(393), I5 =>  inp_feat(456)); 
C_16_S_1_L_5_inst : LUT6 generic map(INIT => "0010001000000000010000001101000010100011011001101100000011010100") port map( O =>C_16_S_1_L_5_out, I0 =>  inp_feat(108), I1 =>  inp_feat(452), I2 =>  inp_feat(20), I3 =>  inp_feat(445), I4 =>  inp_feat(393), I5 =>  inp_feat(456)); 
C_16_S_2_L_0_inst : LUT6 generic map(INIT => "0001100110001000101111110001001110110111000101010111111110100111") port map( O =>C_16_S_2_L_0_out, I0 =>  inp_feat(334), I1 =>  inp_feat(215), I2 =>  inp_feat(352), I3 =>  inp_feat(261), I4 =>  inp_feat(121), I5 =>  inp_feat(485)); 
C_16_S_2_L_1_inst : LUT6 generic map(INIT => "0110101000111111010011000000000010010011111111111100111000001000") port map( O =>C_16_S_2_L_1_out, I0 =>  inp_feat(388), I1 =>  inp_feat(420), I2 =>  inp_feat(445), I3 =>  inp_feat(225), I4 =>  inp_feat(279), I5 =>  inp_feat(263)); 
C_16_S_2_L_2_inst : LUT6 generic map(INIT => "0010110001011101101000110010001011101110111000101010101100001010") port map( O =>C_16_S_2_L_2_out, I0 =>  inp_feat(324), I1 =>  inp_feat(215), I2 =>  inp_feat(244), I3 =>  inp_feat(67), I4 =>  inp_feat(149), I5 =>  inp_feat(190)); 
C_16_S_2_L_3_inst : LUT6 generic map(INIT => "1000010101010011010111110101011100010000000100010000011100111111") port map( O =>C_16_S_2_L_3_out, I0 =>  inp_feat(215), I1 =>  inp_feat(186), I2 =>  inp_feat(199), I3 =>  inp_feat(485), I4 =>  inp_feat(417), I5 =>  inp_feat(430)); 
C_16_S_2_L_4_inst : LUT6 generic map(INIT => "0101110100000011110100010100000011110011000100001110110010000000") port map( O =>C_16_S_2_L_4_out, I0 =>  inp_feat(205), I1 =>  inp_feat(452), I2 =>  inp_feat(137), I3 =>  inp_feat(372), I4 =>  inp_feat(199), I5 =>  inp_feat(417)); 
C_16_S_2_L_5_inst : LUT6 generic map(INIT => "1111000001010111101101100000110100000000001101001001001100000000") port map( O =>C_16_S_2_L_5_out, I0 =>  inp_feat(263), I1 =>  inp_feat(500), I2 =>  inp_feat(332), I3 =>  inp_feat(328), I4 =>  inp_feat(458), I5 =>  inp_feat(17)); 
C_16_S_3_L_0_inst : LUT6 generic map(INIT => "0110000100010101101010100110100001010011001000101010101100001010") port map( O =>C_16_S_3_L_0_out, I0 =>  inp_feat(273), I1 =>  inp_feat(215), I2 =>  inp_feat(244), I3 =>  inp_feat(67), I4 =>  inp_feat(190), I5 =>  inp_feat(149)); 
C_16_S_3_L_1_inst : LUT6 generic map(INIT => "0000101001010100111110110000010011100000000010001111110100000000") port map( O =>C_16_S_3_L_1_out, I0 =>  inp_feat(344), I1 =>  inp_feat(70), I2 =>  inp_feat(224), I3 =>  inp_feat(66), I4 =>  inp_feat(445), I5 =>  inp_feat(395)); 
C_16_S_3_L_2_inst : LUT6 generic map(INIT => "1001001010110001100101001111011111110001010100111111000111110111") port map( O =>C_16_S_3_L_2_out, I0 =>  inp_feat(445), I1 =>  inp_feat(186), I2 =>  inp_feat(363), I3 =>  inp_feat(403), I4 =>  inp_feat(352), I5 =>  inp_feat(226)); 
C_16_S_3_L_3_inst : LUT6 generic map(INIT => "1110100000101010011000001010010000000000000000000000000000110000") port map( O =>C_16_S_3_L_3_out, I0 =>  inp_feat(183), I1 =>  inp_feat(205), I2 =>  inp_feat(62), I3 =>  inp_feat(374), I4 =>  inp_feat(52), I5 =>  inp_feat(405)); 
C_16_S_3_L_4_inst : LUT6 generic map(INIT => "0000000000000100100111100000000010010010000100011110111011001000") port map( O =>C_16_S_3_L_4_out, I0 =>  inp_feat(363), I1 =>  inp_feat(378), I2 =>  inp_feat(81), I3 =>  inp_feat(387), I4 =>  inp_feat(352), I5 =>  inp_feat(403)); 
C_16_S_3_L_5_inst : LUT6 generic map(INIT => "1111001000101101100111011111111100010100000011100000110101001101") port map( O =>C_16_S_3_L_5_out, I0 =>  inp_feat(445), I1 =>  inp_feat(454), I2 =>  inp_feat(186), I3 =>  inp_feat(199), I4 =>  inp_feat(417), I5 =>  inp_feat(430)); 
C_16_S_4_L_0_inst : LUT6 generic map(INIT => "1011010101101011100100111111111100000101000001010000011101111111") port map( O =>C_16_S_4_L_0_out, I0 =>  inp_feat(215), I1 =>  inp_feat(445), I2 =>  inp_feat(186), I3 =>  inp_feat(199), I4 =>  inp_feat(417), I5 =>  inp_feat(430)); 
C_16_S_4_L_1_inst : LUT6 generic map(INIT => "0001010100110111000000110001111110010111011111110001011000010111") port map( O =>C_16_S_4_L_1_out, I0 =>  inp_feat(431), I1 =>  inp_feat(393), I2 =>  inp_feat(353), I3 =>  inp_feat(321), I4 =>  inp_feat(261), I5 =>  inp_feat(111)); 
C_16_S_4_L_2_inst : LUT6 generic map(INIT => "1100101010000001111000110000111000000000000000001010010000000000") port map( O =>C_16_S_4_L_2_out, I0 =>  inp_feat(140), I1 =>  inp_feat(141), I2 =>  inp_feat(50), I3 =>  inp_feat(356), I4 =>  inp_feat(190), I5 =>  inp_feat(442)); 
C_16_S_4_L_3_inst : LUT6 generic map(INIT => "0100000110000000010000001110110010100000000000010100000011000100") port map( O =>C_16_S_4_L_3_out, I0 =>  inp_feat(489), I1 =>  inp_feat(93), I2 =>  inp_feat(299), I3 =>  inp_feat(445), I4 =>  inp_feat(227), I5 =>  inp_feat(281)); 
C_16_S_4_L_4_inst : LUT6 generic map(INIT => "1001000011010001111010110000001000000011110000000000000000000100") port map( O =>C_16_S_4_L_4_out, I0 =>  inp_feat(43), I1 =>  inp_feat(136), I2 =>  inp_feat(324), I3 =>  inp_feat(239), I4 =>  inp_feat(453), I5 =>  inp_feat(430)); 
C_16_S_4_L_5_inst : LUT6 generic map(INIT => "0001011100010111000000001011000011111111000000110000000000000000") port map( O =>C_16_S_4_L_5_out, I0 =>  inp_feat(216), I1 =>  inp_feat(509), I2 =>  inp_feat(145), I3 =>  inp_feat(439), I4 =>  inp_feat(284), I5 =>  inp_feat(460)); 
C_16_S_5_L_0_inst : LUT6 generic map(INIT => "1010100000111111101110001111100100000000000010011100100000000000") port map( O =>C_16_S_5_L_0_out, I0 =>  inp_feat(221), I1 =>  inp_feat(272), I2 =>  inp_feat(107), I3 =>  inp_feat(76), I4 =>  inp_feat(485), I5 =>  inp_feat(430)); 
C_16_S_5_L_1_inst : LUT6 generic map(INIT => "0110001101000111110111110111111100000001000001110000101111111111") port map( O =>C_16_S_5_L_1_out, I0 =>  inp_feat(91), I1 =>  inp_feat(123), I2 =>  inp_feat(215), I3 =>  inp_feat(403), I4 =>  inp_feat(190), I5 =>  inp_feat(442)); 
C_16_S_5_L_2_inst : LUT6 generic map(INIT => "0010101000001010110100101001101010100000111110001010000011110010") port map( O =>C_16_S_5_L_2_out, I0 =>  inp_feat(313), I1 =>  inp_feat(238), I2 =>  inp_feat(231), I3 =>  inp_feat(105), I4 =>  inp_feat(166), I5 =>  inp_feat(474)); 
C_16_S_5_L_3_inst : LUT6 generic map(INIT => "1000100011010000100001000000010010101111000011001001010000000000") port map( O =>C_16_S_5_L_3_out, I0 =>  inp_feat(74), I1 =>  inp_feat(363), I2 =>  inp_feat(447), I3 =>  inp_feat(178), I4 =>  inp_feat(318), I5 =>  inp_feat(344)); 
C_16_S_5_L_4_inst : LUT6 generic map(INIT => "1010001101100111010110110111111100010001000000100000001000010001") port map( O =>C_16_S_5_L_4_out, I0 =>  inp_feat(431), I1 =>  inp_feat(123), I2 =>  inp_feat(194), I3 =>  inp_feat(244), I4 =>  inp_feat(103), I5 =>  inp_feat(479)); 
C_16_S_5_L_5_inst : LUT6 generic map(INIT => "0010000110010000000101000000000100000010010000001111110100000000") port map( O =>C_16_S_5_L_5_out, I0 =>  inp_feat(474), I1 =>  inp_feat(341), I2 =>  inp_feat(56), I3 =>  inp_feat(19), I4 =>  inp_feat(143), I5 =>  inp_feat(295)); 
C_17_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111011001110000011111010100000001000000000000000") port map( O =>C_17_S_0_L_0_out, I0 =>  inp_feat(194), I1 =>  inp_feat(306), I2 =>  inp_feat(392), I3 =>  inp_feat(108), I4 =>  inp_feat(248), I5 =>  inp_feat(239)); 
C_17_S_0_L_1_inst : LUT6 generic map(INIT => "1010100001011110000000001111101000100000001111000000000011000000") port map( O =>C_17_S_0_L_1_out, I0 =>  inp_feat(199), I1 =>  inp_feat(392), I2 =>  inp_feat(186), I3 =>  inp_feat(378), I4 =>  inp_feat(149), I5 =>  inp_feat(497)); 
C_17_S_0_L_2_inst : LUT6 generic map(INIT => "1110001011111101110100110000110001111010000011110000011100000011") port map( O =>C_17_S_0_L_2_out, I0 =>  inp_feat(105), I1 =>  inp_feat(59), I2 =>  inp_feat(420), I3 =>  inp_feat(431), I4 =>  inp_feat(215), I5 =>  inp_feat(353)); 
C_17_S_0_L_3_inst : LUT6 generic map(INIT => "0011011100110010101111011111101000010001001101010011110111111101") port map( O =>C_17_S_0_L_3_out, I0 =>  inp_feat(17), I1 =>  inp_feat(378), I2 =>  inp_feat(277), I3 =>  inp_feat(482), I4 =>  inp_feat(312), I5 =>  inp_feat(241)); 
C_17_S_0_L_4_inst : LUT6 generic map(INIT => "0001101101001000010101010101110110111011001111111111110110011101") port map( O =>C_17_S_0_L_4_out, I0 =>  inp_feat(165), I1 =>  inp_feat(279), I2 =>  inp_feat(427), I3 =>  inp_feat(403), I4 =>  inp_feat(389), I5 =>  inp_feat(415)); 
C_17_S_0_L_5_inst : LUT6 generic map(INIT => "1111111110101001101011110010100010000100000011000000100000001100") port map( O =>C_17_S_0_L_5_out, I0 =>  inp_feat(306), I1 =>  inp_feat(239), I2 =>  inp_feat(48), I3 =>  inp_feat(403), I4 =>  inp_feat(108), I5 =>  inp_feat(241)); 
C_17_S_1_L_0_inst : LUT6 generic map(INIT => "1010100001011110000000001111101000100000001111000000000011000000") port map( O =>C_17_S_1_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(392), I2 =>  inp_feat(186), I3 =>  inp_feat(378), I4 =>  inp_feat(149), I5 =>  inp_feat(497)); 
C_17_S_1_L_1_inst : LUT6 generic map(INIT => "1110001011111101110100110000110001111010000011110000011100000011") port map( O =>C_17_S_1_L_1_out, I0 =>  inp_feat(105), I1 =>  inp_feat(59), I2 =>  inp_feat(420), I3 =>  inp_feat(431), I4 =>  inp_feat(215), I5 =>  inp_feat(353)); 
C_17_S_1_L_2_inst : LUT6 generic map(INIT => "0011011100110010101111011111101000010001001101010011110111111101") port map( O =>C_17_S_1_L_2_out, I0 =>  inp_feat(17), I1 =>  inp_feat(378), I2 =>  inp_feat(277), I3 =>  inp_feat(482), I4 =>  inp_feat(312), I5 =>  inp_feat(241)); 
C_17_S_1_L_3_inst : LUT6 generic map(INIT => "0001101101001000010101010101110110111011001111111111110110011101") port map( O =>C_17_S_1_L_3_out, I0 =>  inp_feat(165), I1 =>  inp_feat(279), I2 =>  inp_feat(427), I3 =>  inp_feat(403), I4 =>  inp_feat(389), I5 =>  inp_feat(415)); 
C_17_S_1_L_4_inst : LUT6 generic map(INIT => "1111111110101001101011110010100010000100000011000000100000001100") port map( O =>C_17_S_1_L_4_out, I0 =>  inp_feat(306), I1 =>  inp_feat(239), I2 =>  inp_feat(48), I3 =>  inp_feat(403), I4 =>  inp_feat(108), I5 =>  inp_feat(241)); 
C_17_S_1_L_5_inst : LUT6 generic map(INIT => "0101001100010010011100100010001011111111101111111111101101101000") port map( O =>C_17_S_1_L_5_out, I0 =>  inp_feat(248), I1 =>  inp_feat(45), I2 =>  inp_feat(121), I3 =>  inp_feat(417), I4 =>  inp_feat(334), I5 =>  inp_feat(419)); 
C_17_S_2_L_0_inst : LUT6 generic map(INIT => "1110001011111011111001110100110110101110010111010000111100000111") port map( O =>C_17_S_2_L_0_out, I0 =>  inp_feat(420), I1 =>  inp_feat(105), I2 =>  inp_feat(402), I3 =>  inp_feat(431), I4 =>  inp_feat(215), I5 =>  inp_feat(353)); 
C_17_S_2_L_1_inst : LUT6 generic map(INIT => "0001110100111111010110101101100000011100111100000100100000000000") port map( O =>C_17_S_2_L_1_out, I0 =>  inp_feat(257), I1 =>  inp_feat(248), I2 =>  inp_feat(169), I3 =>  inp_feat(57), I4 =>  inp_feat(103), I5 =>  inp_feat(7)); 
C_17_S_2_L_2_inst : LUT6 generic map(INIT => "0011110000111101011011001111010111111111111111001111111110011110") port map( O =>C_17_S_2_L_2_out, I0 =>  inp_feat(445), I1 =>  inp_feat(453), I2 =>  inp_feat(406), I3 =>  inp_feat(212), I4 =>  inp_feat(421), I5 =>  inp_feat(208)); 
C_17_S_2_L_3_inst : LUT6 generic map(INIT => "1111101111101111101001111111000101100011111100110101000101010000") port map( O =>C_17_S_2_L_3_out, I0 =>  inp_feat(356), I1 =>  inp_feat(169), I2 =>  inp_feat(103), I3 =>  inp_feat(28), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_17_S_2_L_4_inst : LUT6 generic map(INIT => "0000010010011101001011111111101111110111111111110110111111111111") port map( O =>C_17_S_2_L_4_out, I0 =>  inp_feat(190), I1 =>  inp_feat(294), I2 =>  inp_feat(379), I3 =>  inp_feat(165), I4 =>  inp_feat(248), I5 =>  inp_feat(191)); 
C_17_S_2_L_5_inst : LUT6 generic map(INIT => "1111101010100000101100001010100000100010010110001111100010000000") port map( O =>C_17_S_2_L_5_out, I0 =>  inp_feat(403), I1 =>  inp_feat(392), I2 =>  inp_feat(186), I3 =>  inp_feat(125), I4 =>  inp_feat(263), I5 =>  inp_feat(90)); 
C_17_S_3_L_0_inst : LUT6 generic map(INIT => "1111001011011111110111010001110010111010000001110000111100000001") port map( O =>C_17_S_3_L_0_out, I0 =>  inp_feat(465), I1 =>  inp_feat(59), I2 =>  inp_feat(420), I3 =>  inp_feat(215), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_17_S_3_L_1_inst : LUT6 generic map(INIT => "1010101010100101010010001111100001000000111110001000000010010000") port map( O =>C_17_S_3_L_1_out, I0 =>  inp_feat(334), I1 =>  inp_feat(248), I2 =>  inp_feat(215), I3 =>  inp_feat(14), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_17_S_3_L_2_inst : LUT6 generic map(INIT => "0101100100011111001101111010111001000011111111111110001110101011") port map( O =>C_17_S_3_L_2_out, I0 =>  inp_feat(142), I1 =>  inp_feat(298), I2 =>  inp_feat(217), I3 =>  inp_feat(320), I4 =>  inp_feat(458), I5 =>  inp_feat(229)); 
C_17_S_3_L_3_inst : LUT6 generic map(INIT => "0100000010101000010011001110110011101010011010001111100010101000") port map( O =>C_17_S_3_L_3_out, I0 =>  inp_feat(186), I1 =>  inp_feat(121), I2 =>  inp_feat(199), I3 =>  inp_feat(385), I4 =>  inp_feat(14), I5 =>  inp_feat(502)); 
C_17_S_3_L_4_inst : LUT6 generic map(INIT => "1111101111011101110111111111010100010001110111110100000011110000") port map( O =>C_17_S_3_L_4_out, I0 =>  inp_feat(98), I1 =>  inp_feat(489), I2 =>  inp_feat(218), I3 =>  inp_feat(57), I4 =>  inp_feat(215), I5 =>  inp_feat(186)); 
C_17_S_3_L_5_inst : LUT6 generic map(INIT => "0011101111011111000111111111110100011001110110111111111111111011") port map( O =>C_17_S_3_L_5_out, I0 =>  inp_feat(274), I1 =>  inp_feat(292), I2 =>  inp_feat(359), I3 =>  inp_feat(499), I4 =>  inp_feat(27), I5 =>  inp_feat(232)); 
C_17_S_4_L_0_inst : LUT6 generic map(INIT => "0111111111111010111100111100000001110110101010000001000010000000") port map( O =>C_17_S_4_L_0_out, I0 =>  inp_feat(136), I1 =>  inp_feat(257), I2 =>  inp_feat(352), I3 =>  inp_feat(275), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_17_S_4_L_1_inst : LUT6 generic map(INIT => "0110111111001100100010100000101010101111101001001000110000000000") port map( O =>C_17_S_4_L_1_out, I0 =>  inp_feat(353), I1 =>  inp_feat(403), I2 =>  inp_feat(183), I3 =>  inp_feat(334), I4 =>  inp_feat(215), I5 =>  inp_feat(211)); 
C_17_S_4_L_2_inst : LUT6 generic map(INIT => "0011011000010111111010110011100110111111111111011001001111110010") port map( O =>C_17_S_4_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(175), I2 =>  inp_feat(278), I3 =>  inp_feat(108), I4 =>  inp_feat(229), I5 =>  inp_feat(106)); 
C_17_S_4_L_3_inst : LUT6 generic map(INIT => "1111110111111011111011111111110111111111110000110000000011111111") port map( O =>C_17_S_4_L_3_out, I0 =>  inp_feat(180), I1 =>  inp_feat(204), I2 =>  inp_feat(288), I3 =>  inp_feat(356), I4 =>  inp_feat(431), I5 =>  inp_feat(353)); 
C_17_S_4_L_4_inst : LUT6 generic map(INIT => "1011111101101111111110100001111101011100010101111111111111001111") port map( O =>C_17_S_4_L_4_out, I0 =>  inp_feat(419), I1 =>  inp_feat(405), I2 =>  inp_feat(499), I3 =>  inp_feat(44), I4 =>  inp_feat(37), I5 =>  inp_feat(237)); 
C_17_S_4_L_5_inst : LUT6 generic map(INIT => "0101011101011001000111100101101100000011101111111001101111111010") port map( O =>C_17_S_4_L_5_out, I0 =>  inp_feat(86), I1 =>  inp_feat(279), I2 =>  inp_feat(142), I3 =>  inp_feat(320), I4 =>  inp_feat(458), I5 =>  inp_feat(229)); 
C_17_S_5_L_0_inst : LUT6 generic map(INIT => "0011111101110110111111110001111011111110110111011111110000111110") port map( O =>C_17_S_5_L_0_out, I0 =>  inp_feat(296), I1 =>  inp_feat(475), I2 =>  inp_feat(164), I3 =>  inp_feat(132), I4 =>  inp_feat(285), I5 =>  inp_feat(367)); 
C_17_S_5_L_1_inst : LUT6 generic map(INIT => "1111111011111110011101110110111101111110100000000100011000000000") port map( O =>C_17_S_5_L_1_out, I0 =>  inp_feat(74), I1 =>  inp_feat(303), I2 =>  inp_feat(65), I3 =>  inp_feat(97), I4 =>  inp_feat(215), I5 =>  inp_feat(186)); 
C_17_S_5_L_2_inst : LUT6 generic map(INIT => "1110011001101010111110000010000000001001100010001111100000010010") port map( O =>C_17_S_5_L_2_out, I0 =>  inp_feat(73), I1 =>  inp_feat(288), I2 =>  inp_feat(416), I3 =>  inp_feat(347), I4 =>  inp_feat(295), I5 =>  inp_feat(384)); 
C_17_S_5_L_3_inst : LUT6 generic map(INIT => "0000111000101110010011010010100011011111111111000001111111111110") port map( O =>C_17_S_5_L_3_out, I0 =>  inp_feat(171), I1 =>  inp_feat(338), I2 =>  inp_feat(6), I3 =>  inp_feat(456), I4 =>  inp_feat(237), I5 =>  inp_feat(145)); 
C_17_S_5_L_4_inst : LUT6 generic map(INIT => "1101111011111111011000101101111111101111111011111111001111111111") port map( O =>C_17_S_5_L_4_out, I0 =>  inp_feat(377), I1 =>  inp_feat(480), I2 =>  inp_feat(412), I3 =>  inp_feat(89), I4 =>  inp_feat(35), I5 =>  inp_feat(198)); 
C_17_S_5_L_5_inst : LUT6 generic map(INIT => "1110011100101111011110111000110101010011111111111110001110100011") port map( O =>C_17_S_5_L_5_out, I0 =>  inp_feat(330), I1 =>  inp_feat(298), I2 =>  inp_feat(217), I3 =>  inp_feat(320), I4 =>  inp_feat(458), I5 =>  inp_feat(229)); 
C_18_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000010111000000010101011100000001001101110001011101111111") port map( O =>C_18_S_0_L_0_out, I0 =>  inp_feat(350), I1 =>  inp_feat(83), I2 =>  inp_feat(399), I3 =>  inp_feat(324), I4 =>  inp_feat(373), I5 =>  inp_feat(185)); 
C_18_S_0_L_1_inst : LUT6 generic map(INIT => "0000011101010111010111111111111111110111111111111111111111111111") port map( O =>C_18_S_0_L_1_out, I0 =>  inp_feat(288), I1 =>  inp_feat(449), I2 =>  inp_feat(65), I3 =>  inp_feat(210), I4 =>  inp_feat(26), I5 =>  inp_feat(497)); 
C_18_S_0_L_2_inst : LUT6 generic map(INIT => "0000111001100000110011000000100011111100000000001110110100000100") port map( O =>C_18_S_0_L_2_out, I0 =>  inp_feat(214), I1 =>  inp_feat(456), I2 =>  inp_feat(450), I3 =>  inp_feat(463), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_18_S_0_L_3_inst : LUT6 generic map(INIT => "1111111010111011010110101011111000000010001000100000001010100010") port map( O =>C_18_S_0_L_3_out, I0 =>  inp_feat(137), I1 =>  inp_feat(449), I2 =>  inp_feat(450), I3 =>  inp_feat(404), I4 =>  inp_feat(63), I5 =>  inp_feat(421)); 
C_18_S_0_L_4_inst : LUT6 generic map(INIT => "0010011100000000011011110000000011011111001000011111111100010001") port map( O =>C_18_S_0_L_4_out, I0 =>  inp_feat(26), I1 =>  inp_feat(96), I2 =>  inp_feat(449), I3 =>  inp_feat(84), I4 =>  inp_feat(280), I5 =>  inp_feat(318)); 
C_18_S_0_L_5_inst : LUT6 generic map(INIT => "0101011111011101010001010101110110111111000000000000000000000010") port map( O =>C_18_S_0_L_5_out, I0 =>  inp_feat(328), I1 =>  inp_feat(25), I2 =>  inp_feat(303), I3 =>  inp_feat(260), I4 =>  inp_feat(172), I5 =>  inp_feat(437)); 
C_18_S_1_L_0_inst : LUT6 generic map(INIT => "0000011101010111010111111111111111110111111111111111111111111111") port map( O =>C_18_S_1_L_0_out, I0 =>  inp_feat(288), I1 =>  inp_feat(449), I2 =>  inp_feat(65), I3 =>  inp_feat(210), I4 =>  inp_feat(26), I5 =>  inp_feat(497)); 
C_18_S_1_L_1_inst : LUT6 generic map(INIT => "0000111001100000110011000000100011111100000000001110110100000100") port map( O =>C_18_S_1_L_1_out, I0 =>  inp_feat(214), I1 =>  inp_feat(456), I2 =>  inp_feat(450), I3 =>  inp_feat(463), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_18_S_1_L_2_inst : LUT6 generic map(INIT => "1111111010111011010110101011111000000010001000100000001010100010") port map( O =>C_18_S_1_L_2_out, I0 =>  inp_feat(137), I1 =>  inp_feat(449), I2 =>  inp_feat(450), I3 =>  inp_feat(404), I4 =>  inp_feat(63), I5 =>  inp_feat(421)); 
C_18_S_1_L_3_inst : LUT6 generic map(INIT => "0010011100000000011011110000000011011111001000011111111100010001") port map( O =>C_18_S_1_L_3_out, I0 =>  inp_feat(26), I1 =>  inp_feat(96), I2 =>  inp_feat(449), I3 =>  inp_feat(84), I4 =>  inp_feat(280), I5 =>  inp_feat(318)); 
C_18_S_1_L_4_inst : LUT6 generic map(INIT => "0101011111011101010001010101110110111111000000000000000000000010") port map( O =>C_18_S_1_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(25), I2 =>  inp_feat(303), I3 =>  inp_feat(260), I4 =>  inp_feat(172), I5 =>  inp_feat(437)); 
C_18_S_1_L_5_inst : LUT6 generic map(INIT => "1101010111110011111011001110000000100100110001001000110000000000") port map( O =>C_18_S_1_L_5_out, I0 =>  inp_feat(320), I1 =>  inp_feat(387), I2 =>  inp_feat(363), I3 =>  inp_feat(366), I4 =>  inp_feat(63), I5 =>  inp_feat(46)); 
C_18_S_2_L_0_inst : LUT6 generic map(INIT => "0000010010100100010111000000100111001101000001001100110001001100") port map( O =>C_18_S_2_L_0_out, I0 =>  inp_feat(449), I1 =>  inp_feat(51), I2 =>  inp_feat(289), I3 =>  inp_feat(137), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_18_S_2_L_1_inst : LUT6 generic map(INIT => "1000101001000000011110010000000011110011000100111011101000110000") port map( O =>C_18_S_2_L_1_out, I0 =>  inp_feat(435), I1 =>  inp_feat(318), I2 =>  inp_feat(248), I3 =>  inp_feat(276), I4 =>  inp_feat(280), I5 =>  inp_feat(412)); 
C_18_S_2_L_2_inst : LUT6 generic map(INIT => "0011001110000010110111010001000001111111101001011111111100010111") port map( O =>C_18_S_2_L_2_out, I0 =>  inp_feat(497), I1 =>  inp_feat(412), I2 =>  inp_feat(93), I3 =>  inp_feat(276), I4 =>  inp_feat(136), I5 =>  inp_feat(112)); 
C_18_S_2_L_3_inst : LUT6 generic map(INIT => "0100110111011001110011001100101100001000000001000000000010000001") port map( O =>C_18_S_2_L_3_out, I0 =>  inp_feat(74), I1 =>  inp_feat(50), I2 =>  inp_feat(303), I3 =>  inp_feat(54), I4 =>  inp_feat(486), I5 =>  inp_feat(195)); 
C_18_S_2_L_4_inst : LUT6 generic map(INIT => "0101001101010111010101110010011111000000100001001100100000010001") port map( O =>C_18_S_2_L_4_out, I0 =>  inp_feat(489), I1 =>  inp_feat(303), I2 =>  inp_feat(280), I3 =>  inp_feat(324), I4 =>  inp_feat(83), I5 =>  inp_feat(28)); 
C_18_S_2_L_5_inst : LUT6 generic map(INIT => "1111111101000001111100110111110100010010000000000110010000000010") port map( O =>C_18_S_2_L_5_out, I0 =>  inp_feat(328), I1 =>  inp_feat(126), I2 =>  inp_feat(309), I3 =>  inp_feat(483), I4 =>  inp_feat(399), I5 =>  inp_feat(471)); 
C_18_S_3_L_0_inst : LUT6 generic map(INIT => "0000000100001100011100000100000000010011000011001111001100100000") port map( O =>C_18_S_3_L_0_out, I0 =>  inp_feat(13), I1 =>  inp_feat(115), I2 =>  inp_feat(253), I3 =>  inp_feat(237), I4 =>  inp_feat(361), I5 =>  inp_feat(112)); 
C_18_S_3_L_1_inst : LUT6 generic map(INIT => "0001001111110111110011000110001111011111011101110000000000010001") port map( O =>C_18_S_3_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(489), I2 =>  inp_feat(83), I3 =>  inp_feat(305), I4 =>  inp_feat(246), I5 =>  inp_feat(399)); 
C_18_S_3_L_2_inst : LUT6 generic map(INIT => "1010101000000000100100111100000010110011000010001111011100000000") port map( O =>C_18_S_3_L_2_out, I0 =>  inp_feat(280), I1 =>  inp_feat(328), I2 =>  inp_feat(184), I3 =>  inp_feat(223), I4 =>  inp_feat(210), I5 =>  inp_feat(26)); 
C_18_S_3_L_3_inst : LUT6 generic map(INIT => "0001111101111101000100101111000111111101100101011101000011110000") port map( O =>C_18_S_3_L_3_out, I0 =>  inp_feat(303), I1 =>  inp_feat(502), I2 =>  inp_feat(317), I3 =>  inp_feat(35), I4 =>  inp_feat(65), I5 =>  inp_feat(95)); 
C_18_S_3_L_4_inst : LUT6 generic map(INIT => "0010110001100000110010010000000010001011000000011010111111111001") port map( O =>C_18_S_3_L_4_out, I0 =>  inp_feat(488), I1 =>  inp_feat(279), I2 =>  inp_feat(21), I3 =>  inp_feat(335), I4 =>  inp_feat(196), I5 =>  inp_feat(359)); 
C_18_S_3_L_5_inst : LUT6 generic map(INIT => "1111011101001000000100011100010000000111000000000000100011000000") port map( O =>C_18_S_3_L_5_out, I0 =>  inp_feat(61), I1 =>  inp_feat(214), I2 =>  inp_feat(372), I3 =>  inp_feat(344), I4 =>  inp_feat(389), I5 =>  inp_feat(334)); 
C_18_S_4_L_0_inst : LUT6 generic map(INIT => "0000000001000000111111000100000011011000000100011101110011000100") port map( O =>C_18_S_4_L_0_out, I0 =>  inp_feat(13), I1 =>  inp_feat(363), I2 =>  inp_feat(248), I3 =>  inp_feat(276), I4 =>  inp_feat(280), I5 =>  inp_feat(412)); 
C_18_S_4_L_1_inst : LUT6 generic map(INIT => "1010010001000101110111110010111100000000000000001101110000000100") port map( O =>C_18_S_4_L_1_out, I0 =>  inp_feat(93), I1 =>  inp_feat(418), I2 =>  inp_feat(210), I3 =>  inp_feat(147), I4 =>  inp_feat(13), I5 =>  inp_feat(439)); 
C_18_S_4_L_2_inst : LUT6 generic map(INIT => "0011000000110000101101100001101100100000000000001011000100000000") port map( O =>C_18_S_4_L_2_out, I0 =>  inp_feat(111), I1 =>  inp_feat(25), I2 =>  inp_feat(59), I3 =>  inp_feat(483), I4 =>  inp_feat(229), I5 =>  inp_feat(471)); 
C_18_S_4_L_3_inst : LUT6 generic map(INIT => "0010001001001100110100110000110011110101010110101111011100000000") port map( O =>C_18_S_4_L_3_out, I0 =>  inp_feat(83), I1 =>  inp_feat(350), I2 =>  inp_feat(159), I3 =>  inp_feat(230), I4 =>  inp_feat(299), I5 =>  inp_feat(112)); 
C_18_S_4_L_4_inst : LUT6 generic map(INIT => "1111101000000000100110010000110000000000000000000000000000000010") port map( O =>C_18_S_4_L_4_out, I0 =>  inp_feat(292), I1 =>  inp_feat(479), I2 =>  inp_feat(122), I3 =>  inp_feat(36), I4 =>  inp_feat(483), I5 =>  inp_feat(471)); 
C_18_S_4_L_5_inst : LUT6 generic map(INIT => "0011111100010011000100010000000011101101000001100000000000000100") port map( O =>C_18_S_4_L_5_out, I0 =>  inp_feat(303), I1 =>  inp_feat(136), I2 =>  inp_feat(26), I3 =>  inp_feat(82), I4 =>  inp_feat(172), I5 =>  inp_feat(437)); 
C_18_S_5_L_0_inst : LUT6 generic map(INIT => "0101110001111100110010000110110111101011100000100000000000001000") port map( O =>C_18_S_5_L_0_out, I0 =>  inp_feat(303), I1 =>  inp_feat(246), I2 =>  inp_feat(13), I3 =>  inp_feat(136), I4 =>  inp_feat(60), I5 =>  inp_feat(398)); 
C_18_S_5_L_1_inst : LUT6 generic map(INIT => "1111010111100000000011000000000011110001000000000000000000000000") port map( O =>C_18_S_5_L_1_out, I0 =>  inp_feat(486), I1 =>  inp_feat(124), I2 =>  inp_feat(251), I3 =>  inp_feat(261), I4 =>  inp_feat(50), I5 =>  inp_feat(382)); 
C_18_S_5_L_2_inst : LUT6 generic map(INIT => "0000100111000000010111111101100000000000000010001111001111001010") port map( O =>C_18_S_5_L_2_out, I0 =>  inp_feat(437), I1 =>  inp_feat(130), I2 =>  inp_feat(229), I3 =>  inp_feat(125), I4 =>  inp_feat(244), I5 =>  inp_feat(382)); 
C_18_S_5_L_3_inst : LUT6 generic map(INIT => "1011110011001011100010001010000100000000000001100000000010000001") port map( O =>C_18_S_5_L_3_out, I0 =>  inp_feat(310), I1 =>  inp_feat(116), I2 =>  inp_feat(68), I3 =>  inp_feat(189), I4 =>  inp_feat(74), I5 =>  inp_feat(330)); 
C_18_S_5_L_4_inst : LUT6 generic map(INIT => "0110111101010100111000100000000000010010000010000011000010000000") port map( O =>C_18_S_5_L_4_out, I0 =>  inp_feat(27), I1 =>  inp_feat(77), I2 =>  inp_feat(196), I3 =>  inp_feat(5), I4 =>  inp_feat(205), I5 =>  inp_feat(127)); 
C_18_S_5_L_5_inst : LUT6 generic map(INIT => "0010100010010010000010111100111000000010000000000000000011000000") port map( O =>C_18_S_5_L_5_out, I0 =>  inp_feat(499), I1 =>  inp_feat(458), I2 =>  inp_feat(399), I3 =>  inp_feat(359), I4 =>  inp_feat(196), I5 =>  inp_feat(281)); 
C_19_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000010101000000000000011100000001001111110011011111111111") port map( O =>C_19_S_0_L_0_out, I0 =>  inp_feat(83), I1 =>  inp_feat(318), I2 =>  inp_feat(399), I3 =>  inp_feat(324), I4 =>  inp_feat(373), I5 =>  inp_feat(185)); 
C_19_S_0_L_1_inst : LUT6 generic map(INIT => "0001000011110000100110001111001011110001111100011111000011110010") port map( O =>C_19_S_0_L_1_out, I0 =>  inp_feat(91), I1 =>  inp_feat(328), I2 =>  inp_feat(374), I3 =>  inp_feat(210), I4 =>  inp_feat(65), I5 =>  inp_feat(497)); 
C_19_S_0_L_2_inst : LUT6 generic map(INIT => "1000100000000000000110001100000010001101111100011100100011101100") port map( O =>C_19_S_0_L_2_out, I0 =>  inp_feat(435), I1 =>  inp_feat(434), I2 =>  inp_feat(248), I3 =>  inp_feat(65), I4 =>  inp_feat(210), I5 =>  inp_feat(328)); 
C_19_S_0_L_3_inst : LUT6 generic map(INIT => "0100001101010101111100011111000111111011111111101111000111111111") port map( O =>C_19_S_0_L_3_out, I0 =>  inp_feat(328), I1 =>  inp_feat(399), I2 =>  inp_feat(107), I3 =>  inp_feat(350), I4 =>  inp_feat(280), I5 =>  inp_feat(112)); 
C_19_S_0_L_4_inst : LUT6 generic map(INIT => "0111111101010010010100001100000001110000010000000000000011000000") port map( O =>C_19_S_0_L_4_out, I0 =>  inp_feat(59), I1 =>  inp_feat(83), I2 =>  inp_feat(344), I3 =>  inp_feat(427), I4 =>  inp_feat(11), I5 =>  inp_feat(127)); 
C_19_S_0_L_5_inst : LUT6 generic map(INIT => "1100010001110111101010001101000101000000110011011100000011011100") port map( O =>C_19_S_0_L_5_out, I0 =>  inp_feat(126), I1 =>  inp_feat(245), I2 =>  inp_feat(119), I3 =>  inp_feat(210), I4 =>  inp_feat(361), I5 =>  inp_feat(35)); 
C_19_S_1_L_0_inst : LUT6 generic map(INIT => "0001000011110000100110001111001011110001111100011111000011110010") port map( O =>C_19_S_1_L_0_out, I0 =>  inp_feat(91), I1 =>  inp_feat(328), I2 =>  inp_feat(374), I3 =>  inp_feat(210), I4 =>  inp_feat(65), I5 =>  inp_feat(497)); 
C_19_S_1_L_1_inst : LUT6 generic map(INIT => "1000100000000000000110001100000010001101111100011100100011101100") port map( O =>C_19_S_1_L_1_out, I0 =>  inp_feat(435), I1 =>  inp_feat(434), I2 =>  inp_feat(248), I3 =>  inp_feat(65), I4 =>  inp_feat(210), I5 =>  inp_feat(328)); 
C_19_S_1_L_2_inst : LUT6 generic map(INIT => "0100001101010101111100011111000111111011111111101111000111111111") port map( O =>C_19_S_1_L_2_out, I0 =>  inp_feat(328), I1 =>  inp_feat(399), I2 =>  inp_feat(107), I3 =>  inp_feat(350), I4 =>  inp_feat(280), I5 =>  inp_feat(112)); 
C_19_S_1_L_3_inst : LUT6 generic map(INIT => "0111111101010010010100001100000001110000010000000000000011000000") port map( O =>C_19_S_1_L_3_out, I0 =>  inp_feat(59), I1 =>  inp_feat(83), I2 =>  inp_feat(344), I3 =>  inp_feat(427), I4 =>  inp_feat(11), I5 =>  inp_feat(127)); 
C_19_S_1_L_4_inst : LUT6 generic map(INIT => "1100010001110111101010001101000101000000110011011100000011011100") port map( O =>C_19_S_1_L_4_out, I0 =>  inp_feat(126), I1 =>  inp_feat(245), I2 =>  inp_feat(119), I3 =>  inp_feat(210), I4 =>  inp_feat(361), I5 =>  inp_feat(35)); 
C_19_S_1_L_5_inst : LUT6 generic map(INIT => "0100100111010001000110001101011100000000110001001100000011010100") port map( O =>C_19_S_1_L_5_out, I0 =>  inp_feat(126), I1 =>  inp_feat(4), I2 =>  inp_feat(119), I3 =>  inp_feat(210), I4 =>  inp_feat(361), I5 =>  inp_feat(35)); 
C_19_S_2_L_0_inst : LUT6 generic map(INIT => "1101110101010111001011111111111110101011101101110011011111111111") port map( O =>C_19_S_2_L_0_out, I0 =>  inp_feat(450), I1 =>  inp_feat(489), I2 =>  inp_feat(83), I3 =>  inp_feat(324), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_2_L_1_inst : LUT6 generic map(INIT => "0100000000000010101001001010000011100010101100001010001000100000") port map( O =>C_19_S_2_L_1_out, I0 =>  inp_feat(304), I1 =>  inp_feat(328), I2 =>  inp_feat(482), I3 =>  inp_feat(473), I4 =>  inp_feat(489), I5 =>  inp_feat(350)); 
C_19_S_2_L_2_inst : LUT6 generic map(INIT => "1111010111111011111101110000001001010001000100000010101000000000") port map( O =>C_19_S_2_L_2_out, I0 =>  inp_feat(485), I1 =>  inp_feat(497), I2 =>  inp_feat(266), I3 =>  inp_feat(339), I4 =>  inp_feat(11), I5 =>  inp_feat(127)); 
C_19_S_2_L_3_inst : LUT6 generic map(INIT => "0001110000010011000110010101111101010001010111110001111111111111") port map( O =>C_19_S_2_L_3_out, I0 =>  inp_feat(280), I1 =>  inp_feat(26), I2 =>  inp_feat(318), I3 =>  inp_feat(210), I4 =>  inp_feat(65), I5 =>  inp_feat(35)); 
C_19_S_2_L_4_inst : LUT6 generic map(INIT => "1010101010011000110000011101000011001011110001001100000011001100") port map( O =>C_19_S_2_L_4_out, I0 =>  inp_feat(446), I1 =>  inp_feat(334), I2 =>  inp_feat(180), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_2_L_5_inst : LUT6 generic map(INIT => "0011001100010111010101111011111111100101010111110001110111111111") port map( O =>C_19_S_2_L_5_out, I0 =>  inp_feat(328), I1 =>  inp_feat(445), I2 =>  inp_feat(26), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_3_L_0_inst : LUT6 generic map(INIT => "1111011110110000111100101111000011111001111100001011000011110000") port map( O =>C_19_S_3_L_0_out, I0 =>  inp_feat(214), I1 =>  inp_feat(257), I2 =>  inp_feat(317), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_3_L_1_inst : LUT6 generic map(INIT => "0000011000101011000010111011111000001010111010110010101110111111") port map( O =>C_19_S_3_L_1_out, I0 =>  inp_feat(195), I1 =>  inp_feat(318), I2 =>  inp_feat(65), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_3_L_2_inst : LUT6 generic map(INIT => "1111111011001100110100101100110001011101010001001100000011100110") port map( O =>C_19_S_3_L_2_out, I0 =>  inp_feat(450), I1 =>  inp_feat(275), I2 =>  inp_feat(42), I3 =>  inp_feat(210), I4 =>  inp_feat(13), I5 =>  inp_feat(127)); 
C_19_S_3_L_3_inst : LUT6 generic map(INIT => "1000000110000010000101101101011000000000000001010000000100000010") port map( O =>C_19_S_3_L_3_out, I0 =>  inp_feat(441), I1 =>  inp_feat(439), I2 =>  inp_feat(326), I3 =>  inp_feat(60), I4 =>  inp_feat(234), I5 =>  inp_feat(451)); 
C_19_S_3_L_4_inst : LUT6 generic map(INIT => "0000010000001100010011000001110011011100000101001101110100001100") port map( O =>C_19_S_3_L_4_out, I0 =>  inp_feat(214), I1 =>  inp_feat(456), I2 =>  inp_feat(112), I3 =>  inp_feat(426), I4 =>  inp_feat(303), I5 =>  inp_feat(272)); 
C_19_S_3_L_5_inst : LUT6 generic map(INIT => "1101111111011110010001100001010111000000000001110000000000110000") port map( O =>C_19_S_3_L_5_out, I0 =>  inp_feat(170), I1 =>  inp_feat(461), I2 =>  inp_feat(1), I3 =>  inp_feat(92), I4 =>  inp_feat(344), I5 =>  inp_feat(219)); 
C_19_S_4_L_0_inst : LUT6 generic map(INIT => "1001000000000101000101110111111101010001011111110001111111111111") port map( O =>C_19_S_4_L_0_out, I0 =>  inp_feat(65), I1 =>  inp_feat(257), I2 =>  inp_feat(83), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_4_L_1_inst : LUT6 generic map(INIT => "0010010000101110000110001111010111010010111100101111000011110111") port map( O =>C_19_S_4_L_1_out, I0 =>  inp_feat(168), I1 =>  inp_feat(412), I2 =>  inp_feat(180), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_4_L_2_inst : LUT6 generic map(INIT => "1000101001101011101000101010001000000010000000001100100000000001") port map( O =>C_19_S_4_L_2_out, I0 =>  inp_feat(151), I1 =>  inp_feat(324), I2 =>  inp_feat(143), I3 =>  inp_feat(318), I4 =>  inp_feat(332), I5 =>  inp_feat(292)); 
C_19_S_4_L_3_inst : LUT6 generic map(INIT => "0000100010001000010011000101100010101100100010001100110100001010") port map( O =>C_19_S_4_L_3_out, I0 =>  inp_feat(219), I1 =>  inp_feat(46), I2 =>  inp_feat(95), I3 =>  inp_feat(248), I4 =>  inp_feat(210), I5 =>  inp_feat(303)); 
C_19_S_4_L_4_inst : LUT6 generic map(INIT => "1101010100110111001100011111011100111101000000110001000100110011") port map( O =>C_19_S_4_L_4_out, I0 =>  inp_feat(210), I1 =>  inp_feat(328), I2 =>  inp_feat(35), I3 =>  inp_feat(96), I4 =>  inp_feat(111), I5 =>  inp_feat(266)); 
C_19_S_4_L_5_inst : LUT6 generic map(INIT => "0000101000011001010010100000101111000111000010001110101000000000") port map( O =>C_19_S_4_L_5_out, I0 =>  inp_feat(180), I1 =>  inp_feat(20), I2 =>  inp_feat(60), I3 =>  inp_feat(275), I4 =>  inp_feat(210), I5 =>  inp_feat(328)); 
C_19_S_5_L_0_inst : LUT6 generic map(INIT => "0100000101110111011001111011111110010101010111110011111111111111") port map( O =>C_19_S_5_L_0_out, I0 =>  inp_feat(361), I1 =>  inp_feat(445), I2 =>  inp_feat(26), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_5_L_1_inst : LUT6 generic map(INIT => "1000001011000011110101010111111101010111001111110011111111111111") port map( O =>C_19_S_5_L_1_out, I0 =>  inp_feat(324), I1 =>  inp_feat(445), I2 =>  inp_feat(26), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(35)); 
C_19_S_5_L_2_inst : LUT6 generic map(INIT => "1101100100010010010101000100000011101010011000001111011100000000") port map( O =>C_19_S_5_L_2_out, I0 =>  inp_feat(373), I1 =>  inp_feat(407), I2 =>  inp_feat(191), I3 =>  inp_feat(386), I4 =>  inp_feat(361), I5 =>  inp_feat(83)); 
C_19_S_5_L_3_inst : LUT6 generic map(INIT => "0101001000001101000001001010110001110100000000100000000000000000") port map( O =>C_19_S_5_L_3_out, I0 =>  inp_feat(322), I1 =>  inp_feat(498), I2 =>  inp_feat(440), I3 =>  inp_feat(426), I4 =>  inp_feat(451), I5 =>  inp_feat(234)); 
C_19_S_5_L_4_inst : LUT6 generic map(INIT => "1101000011000101010100100000011000000110110110010000001000000010") port map( O =>C_19_S_5_L_4_out, I0 =>  inp_feat(449), I1 =>  inp_feat(439), I2 =>  inp_feat(326), I3 =>  inp_feat(60), I4 =>  inp_feat(451), I5 =>  inp_feat(234)); 
C_19_S_5_L_5_inst : LUT6 generic map(INIT => "1000111010100000000100001111100100010010100000000000000000000000") port map( O =>C_19_S_5_L_5_out, I0 =>  inp_feat(230), I1 =>  inp_feat(413), I2 =>  inp_feat(263), I3 =>  inp_feat(470), I4 =>  inp_feat(375), I5 =>  inp_feat(304)); 
C_20_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111101010111111111111100011111100110000001100100000000000") port map( O =>C_20_S_0_L_0_out, I0 =>  inp_feat(83), I1 =>  inp_feat(318), I2 =>  inp_feat(399), I3 =>  inp_feat(324), I4 =>  inp_feat(373), I5 =>  inp_feat(185)); 
C_20_S_0_L_1_inst : LUT6 generic map(INIT => "1100100011000100111111101111111100000000010000011110000011101111") port map( O =>C_20_S_0_L_1_out, I0 =>  inp_feat(13), I1 =>  inp_feat(489), I2 =>  inp_feat(318), I3 =>  inp_feat(413), I4 =>  inp_feat(183), I5 =>  inp_feat(35)); 
C_20_S_0_L_2_inst : LUT6 generic map(INIT => "0100000011000100010101001000100011111111111110000111111011001000") port map( O =>C_20_S_0_L_2_out, I0 =>  inp_feat(96), I1 =>  inp_feat(83), I2 =>  inp_feat(65), I3 =>  inp_feat(280), I4 =>  inp_feat(325), I5 =>  inp_feat(183)); 
C_20_S_0_L_3_inst : LUT6 generic map(INIT => "1111101001101010111011101000000000001100111010001000000000000000") port map( O =>C_20_S_0_L_3_out, I0 =>  inp_feat(210), I1 =>  inp_feat(26), I2 =>  inp_feat(328), I3 =>  inp_feat(257), I4 =>  inp_feat(350), I5 =>  inp_feat(280)); 
C_20_S_0_L_4_inst : LUT6 generic map(INIT => "0111000001011110001010001111110010101000011110001000000011101000") port map( O =>C_20_S_0_L_4_out, I0 =>  inp_feat(489), I1 =>  inp_feat(65), I2 =>  inp_feat(83), I3 =>  inp_feat(468), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_20_S_0_L_5_inst : LUT6 generic map(INIT => "1101011101110001011010111100011111101111111111111111111111110111") port map( O =>C_20_S_0_L_5_out, I0 =>  inp_feat(418), I1 =>  inp_feat(74), I2 =>  inp_feat(449), I3 =>  inp_feat(112), I4 =>  inp_feat(59), I5 =>  inp_feat(312)); 
C_20_S_1_L_0_inst : LUT6 generic map(INIT => "1100100011000100111111101111111100000000010000011110000011101111") port map( O =>C_20_S_1_L_0_out, I0 =>  inp_feat(13), I1 =>  inp_feat(489), I2 =>  inp_feat(318), I3 =>  inp_feat(413), I4 =>  inp_feat(183), I5 =>  inp_feat(35)); 
C_20_S_1_L_1_inst : LUT6 generic map(INIT => "0100000011000100010101001000100011111111111110000111111011001000") port map( O =>C_20_S_1_L_1_out, I0 =>  inp_feat(96), I1 =>  inp_feat(83), I2 =>  inp_feat(65), I3 =>  inp_feat(280), I4 =>  inp_feat(325), I5 =>  inp_feat(183)); 
C_20_S_1_L_2_inst : LUT6 generic map(INIT => "1111101001101010111011101000000000001100111010001000000000000000") port map( O =>C_20_S_1_L_2_out, I0 =>  inp_feat(210), I1 =>  inp_feat(26), I2 =>  inp_feat(328), I3 =>  inp_feat(257), I4 =>  inp_feat(350), I5 =>  inp_feat(280)); 
C_20_S_1_L_3_inst : LUT6 generic map(INIT => "0111000001011110001010001111110010101000011110001000000011101000") port map( O =>C_20_S_1_L_3_out, I0 =>  inp_feat(489), I1 =>  inp_feat(65), I2 =>  inp_feat(83), I3 =>  inp_feat(468), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_20_S_1_L_4_inst : LUT6 generic map(INIT => "1101011101110001011010111100011111101111111111111111111111110111") port map( O =>C_20_S_1_L_4_out, I0 =>  inp_feat(418), I1 =>  inp_feat(74), I2 =>  inp_feat(449), I3 =>  inp_feat(112), I4 =>  inp_feat(59), I5 =>  inp_feat(312)); 
C_20_S_1_L_5_inst : LUT6 generic map(INIT => "0010011101100111101010111110001111011001111011111111111111111111") port map( O =>C_20_S_1_L_5_out, I0 =>  inp_feat(203), I1 =>  inp_feat(102), I2 =>  inp_feat(449), I3 =>  inp_feat(112), I4 =>  inp_feat(59), I5 =>  inp_feat(312)); 
C_20_S_2_L_0_inst : LUT6 generic map(INIT => "0111010011000000110010000100000011111010111110001110100010000000") port map( O =>C_20_S_2_L_0_out, I0 =>  inp_feat(280), I1 =>  inp_feat(497), I2 =>  inp_feat(65), I3 =>  inp_feat(210), I4 =>  inp_feat(35), I5 =>  inp_feat(183)); 
C_20_S_2_L_1_inst : LUT6 generic map(INIT => "1110111001001011101100110000001000110010111100101011001100000000") port map( O =>C_20_S_2_L_1_out, I0 =>  inp_feat(361), I1 =>  inp_feat(287), I2 =>  inp_feat(328), I3 =>  inp_feat(324), I4 =>  inp_feat(350), I5 =>  inp_feat(497)); 
C_20_S_2_L_2_inst : LUT6 generic map(INIT => "1010010000101110101011110000111000111111000011000000111000000100") port map( O =>C_20_S_2_L_2_out, I0 =>  inp_feat(210), I1 =>  inp_feat(350), I2 =>  inp_feat(50), I3 =>  inp_feat(280), I4 =>  inp_feat(303), I5 =>  inp_feat(420)); 
C_20_S_2_L_3_inst : LUT6 generic map(INIT => "0101001111110010010100010111000001100010101000101000000000000000") port map( O =>C_20_S_2_L_3_out, I0 =>  inp_feat(185), I1 =>  inp_feat(183), I2 =>  inp_feat(83), I3 =>  inp_feat(324), I4 =>  inp_feat(350), I5 =>  inp_feat(388)); 
C_20_S_2_L_4_inst : LUT6 generic map(INIT => "1101100111110001110101001111111001101100111111000010000011111010") port map( O =>C_20_S_2_L_4_out, I0 =>  inp_feat(432), I1 =>  inp_feat(394), I2 =>  inp_feat(2), I3 =>  inp_feat(473), I4 =>  inp_feat(350), I5 =>  inp_feat(280)); 
C_20_S_2_L_5_inst : LUT6 generic map(INIT => "0011010011001100111111101111111101110000110000001111111111101111") port map( O =>C_20_S_2_L_5_out, I0 =>  inp_feat(104), I1 =>  inp_feat(413), I2 =>  inp_feat(497), I3 =>  inp_feat(101), I4 =>  inp_feat(18), I5 =>  inp_feat(388)); 
C_20_S_3_L_0_inst : LUT6 generic map(INIT => "1111011111100011100011100000111100101100000011000000111000000000") port map( O =>C_20_S_3_L_0_out, I0 =>  inp_feat(210), I1 =>  inp_feat(26), I2 =>  inp_feat(169), I3 =>  inp_feat(324), I4 =>  inp_feat(350), I5 =>  inp_feat(497)); 
C_20_S_3_L_1_inst : LUT6 generic map(INIT => "1101010000110010010011101111011001000000001000000101010010100000") port map( O =>C_20_S_3_L_1_out, I0 =>  inp_feat(206), I1 =>  inp_feat(106), I2 =>  inp_feat(189), I3 =>  inp_feat(237), I4 =>  inp_feat(350), I5 =>  inp_feat(280)); 
C_20_S_3_L_2_inst : LUT6 generic map(INIT => "0100010111110101111011011111110101100100000100001110100000000000") port map( O =>C_20_S_3_L_2_out, I0 =>  inp_feat(419), I1 =>  inp_feat(259), I2 =>  inp_feat(83), I3 =>  inp_feat(185), I4 =>  inp_feat(18), I5 =>  inp_feat(388)); 
C_20_S_3_L_3_inst : LUT6 generic map(INIT => "1100011010101111111001010000100001010000000010100000100000000000") port map( O =>C_20_S_3_L_3_out, I0 =>  inp_feat(328), I1 =>  inp_feat(126), I2 =>  inp_feat(403), I3 =>  inp_feat(280), I4 =>  inp_feat(350), I5 =>  inp_feat(388)); 
C_20_S_3_L_4_inst : LUT6 generic map(INIT => "0000101011001100010001011101110100001010000000000000111111111110") port map( O =>C_20_S_3_L_4_out, I0 =>  inp_feat(117), I1 =>  inp_feat(458), I2 =>  inp_feat(376), I3 =>  inp_feat(8), I4 =>  inp_feat(450), I5 =>  inp_feat(172)); 
C_20_S_3_L_5_inst : LUT6 generic map(INIT => "0011110111111100001111011011101111111111111111110011110111111101") port map( O =>C_20_S_3_L_5_out, I0 =>  inp_feat(374), I1 =>  inp_feat(427), I2 =>  inp_feat(100), I3 =>  inp_feat(307), I4 =>  inp_feat(500), I5 =>  inp_feat(456)); 
C_20_S_4_L_0_inst : LUT6 generic map(INIT => "1011101100001110111101111000111101111011001111110101111111111111") port map( O =>C_20_S_4_L_0_out, I0 =>  inp_feat(394), I1 =>  inp_feat(50), I2 =>  inp_feat(419), I3 =>  inp_feat(386), I4 =>  inp_feat(361), I5 =>  inp_feat(83)); 
C_20_S_4_L_1_inst : LUT6 generic map(INIT => "1111010111101000111000001000000000001100010000001100110011110000") port map( O =>C_20_S_4_L_1_out, I0 =>  inp_feat(83), I1 =>  inp_feat(318), I2 =>  inp_feat(210), I3 =>  inp_feat(65), I4 =>  inp_feat(35), I5 =>  inp_feat(11)); 
C_20_S_4_L_2_inst : LUT6 generic map(INIT => "0010001001111110001000101111111011111111101111110101001000101111") port map( O =>C_20_S_4_L_2_out, I0 =>  inp_feat(115), I1 =>  inp_feat(192), I2 =>  inp_feat(507), I3 =>  inp_feat(165), I4 =>  inp_feat(219), I5 =>  inp_feat(321)); 
C_20_S_4_L_3_inst : LUT6 generic map(INIT => "1010011011110010101110111111001001110000111010100110001111110101") port map( O =>C_20_S_4_L_3_out, I0 =>  inp_feat(418), I1 =>  inp_feat(456), I2 =>  inp_feat(431), I3 =>  inp_feat(230), I4 =>  inp_feat(173), I5 =>  inp_feat(388)); 
C_20_S_4_L_4_inst : LUT6 generic map(INIT => "1110101101011111110111110100111100110010011011111101111110001111") port map( O =>C_20_S_4_L_4_out, I0 =>  inp_feat(488), I1 =>  inp_feat(272), I2 =>  inp_feat(10), I3 =>  inp_feat(210), I4 =>  inp_feat(26), I5 =>  inp_feat(142)); 
C_20_S_4_L_5_inst : LUT6 generic map(INIT => "0101010100011111111111111101101000000000000000101011001111100011") port map( O =>C_20_S_4_L_5_out, I0 =>  inp_feat(59), I1 =>  inp_feat(151), I2 =>  inp_feat(437), I3 =>  inp_feat(377), I4 =>  inp_feat(390), I5 =>  inp_feat(111)); 
C_20_S_5_L_0_inst : LUT6 generic map(INIT => "0111111011111100011010101100000001111100100000000100000000000000") port map( O =>C_20_S_5_L_0_out, I0 =>  inp_feat(303), I1 =>  inp_feat(210), I2 =>  inp_feat(26), I3 =>  inp_feat(373), I4 =>  inp_feat(350), I5 =>  inp_feat(76)); 
C_20_S_5_L_1_inst : LUT6 generic map(INIT => "1011101101111011110101010010000001000010111000000000000010100000") port map( O =>C_20_S_5_L_1_out, I0 =>  inp_feat(304), I1 =>  inp_feat(510), I2 =>  inp_feat(350), I3 =>  inp_feat(166), I4 =>  inp_feat(280), I5 =>  inp_feat(388)); 
C_20_S_5_L_2_inst : LUT6 generic map(INIT => "1010111010100111111101110101001111100100100011100011001111110011") port map( O =>C_20_S_5_L_2_out, I0 =>  inp_feat(105), I1 =>  inp_feat(464), I2 =>  inp_feat(273), I3 =>  inp_feat(335), I4 =>  inp_feat(350), I5 =>  inp_feat(65)); 
C_20_S_5_L_3_inst : LUT6 generic map(INIT => "0011111101011011011111111111111000001010011011010101101101011110") port map( O =>C_20_S_5_L_3_out, I0 =>  inp_feat(173), I1 =>  inp_feat(226), I2 =>  inp_feat(37), I3 =>  inp_feat(307), I4 =>  inp_feat(156), I5 =>  inp_feat(111)); 
C_20_S_5_L_4_inst : LUT6 generic map(INIT => "1101110101111110001010110010111100110100101101110011000110111111") port map( O =>C_20_S_5_L_4_out, I0 =>  inp_feat(63), I1 =>  inp_feat(334), I2 =>  inp_feat(393), I3 =>  inp_feat(26), I4 =>  inp_feat(35), I5 =>  inp_feat(227)); 
C_20_S_5_L_5_inst : LUT6 generic map(INIT => "0010011110001011101000110011000011001111111011101010111100110000") port map( O =>C_20_S_5_L_5_out, I0 =>  inp_feat(172), I1 =>  inp_feat(478), I2 =>  inp_feat(139), I3 =>  inp_feat(330), I4 =>  inp_feat(371), I5 =>  inp_feat(256)); 
C_21_S_0_L_0_inst : LUT6 generic map(INIT => "0000000100010111000101110111111100000001001111110111111101111111") port map( O =>C_21_S_0_L_0_out, I0 =>  inp_feat(280), I1 =>  inp_feat(399), I2 =>  inp_feat(318), I3 =>  inp_feat(324), I4 =>  inp_feat(185), I5 =>  inp_feat(35)); 
C_21_S_0_L_1_inst : LUT6 generic map(INIT => "0000000000001010110100100000000001001010100011100101110000001000") port map( O =>C_21_S_0_L_1_out, I0 =>  inp_feat(248), I1 =>  inp_feat(345), I2 =>  inp_feat(324), I3 =>  inp_feat(350), I4 =>  inp_feat(227), I5 =>  inp_feat(489)); 
C_21_S_0_L_2_inst : LUT6 generic map(INIT => "0000000010000000000100111000000101111111010100011111111111111011") port map( O =>C_21_S_0_L_2_out, I0 =>  inp_feat(26), I1 =>  inp_feat(257), I2 =>  inp_feat(86), I3 =>  inp_feat(321), I4 =>  inp_feat(373), I5 =>  inp_feat(350)); 
C_21_S_0_L_3_inst : LUT6 generic map(INIT => "1010000000000100000001010001110111100100000011010101111111111111") port map( O =>C_21_S_0_L_3_out, I0 =>  inp_feat(35), I1 =>  inp_feat(15), I2 =>  inp_feat(112), I3 =>  inp_feat(449), I4 =>  inp_feat(83), I5 =>  inp_feat(361)); 
C_21_S_0_L_4_inst : LUT6 generic map(INIT => "0000011010000010100000111011101110000100000010111010101110111111") port map( O =>C_21_S_0_L_4_out, I0 =>  inp_feat(173), I1 =>  inp_feat(65), I2 =>  inp_feat(210), I3 =>  inp_feat(112), I4 =>  inp_feat(83), I5 =>  inp_feat(361)); 
C_21_S_0_L_5_inst : LUT6 generic map(INIT => "1000110111100011100010111101111111001001110011110001011101111111") port map( O =>C_21_S_0_L_5_out, I0 =>  inp_feat(324), I1 =>  inp_feat(185), I2 =>  inp_feat(83), I3 =>  inp_feat(373), I4 =>  inp_feat(450), I5 =>  inp_feat(509)); 
C_21_S_1_L_0_inst : LUT6 generic map(INIT => "0000000000001010110100100000000001001010100011100101110000001000") port map( O =>C_21_S_1_L_0_out, I0 =>  inp_feat(248), I1 =>  inp_feat(345), I2 =>  inp_feat(324), I3 =>  inp_feat(350), I4 =>  inp_feat(227), I5 =>  inp_feat(489)); 
C_21_S_1_L_1_inst : LUT6 generic map(INIT => "0000000010000000000100111000000101111111010100011111111111111011") port map( O =>C_21_S_1_L_1_out, I0 =>  inp_feat(26), I1 =>  inp_feat(257), I2 =>  inp_feat(86), I3 =>  inp_feat(321), I4 =>  inp_feat(373), I5 =>  inp_feat(350)); 
C_21_S_1_L_2_inst : LUT6 generic map(INIT => "1010000000000100000001010001110111100100000011010101111111111111") port map( O =>C_21_S_1_L_2_out, I0 =>  inp_feat(35), I1 =>  inp_feat(15), I2 =>  inp_feat(112), I3 =>  inp_feat(449), I4 =>  inp_feat(83), I5 =>  inp_feat(361)); 
C_21_S_1_L_3_inst : LUT6 generic map(INIT => "0000011010000010100000111011101110000100000010111010101110111111") port map( O =>C_21_S_1_L_3_out, I0 =>  inp_feat(173), I1 =>  inp_feat(65), I2 =>  inp_feat(210), I3 =>  inp_feat(112), I4 =>  inp_feat(83), I5 =>  inp_feat(361)); 
C_21_S_1_L_4_inst : LUT6 generic map(INIT => "1000110111100011100010111101111111001001110011110001011101111111") port map( O =>C_21_S_1_L_4_out, I0 =>  inp_feat(324), I1 =>  inp_feat(185), I2 =>  inp_feat(83), I3 =>  inp_feat(373), I4 =>  inp_feat(450), I5 =>  inp_feat(509)); 
C_21_S_1_L_5_inst : LUT6 generic map(INIT => "0000101100010011011000110001011100010001100111110001111101111111") port map( O =>C_21_S_1_L_5_out, I0 =>  inp_feat(210), I1 =>  inp_feat(65), I2 =>  inp_feat(83), I3 =>  inp_feat(303), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_2_L_0_inst : LUT6 generic map(INIT => "0000000010000000000100111000100101111111010100011111111111111011") port map( O =>C_21_S_2_L_0_out, I0 =>  inp_feat(26), I1 =>  inp_feat(257), I2 =>  inp_feat(86), I3 =>  inp_feat(321), I4 =>  inp_feat(373), I5 =>  inp_feat(350)); 
C_21_S_2_L_1_inst : LUT6 generic map(INIT => "1010000000000100000000010001110111100100000011010101111111111111") port map( O =>C_21_S_2_L_1_out, I0 =>  inp_feat(35), I1 =>  inp_feat(15), I2 =>  inp_feat(112), I3 =>  inp_feat(449), I4 =>  inp_feat(83), I5 =>  inp_feat(361)); 
C_21_S_2_L_2_inst : LUT6 generic map(INIT => "0000011010000010100000111011101110000100000010111010101110111111") port map( O =>C_21_S_2_L_2_out, I0 =>  inp_feat(173), I1 =>  inp_feat(65), I2 =>  inp_feat(210), I3 =>  inp_feat(112), I4 =>  inp_feat(83), I5 =>  inp_feat(361)); 
C_21_S_2_L_3_inst : LUT6 generic map(INIT => "0010110011000101111011011100110111101100110011010100110111011101") port map( O =>C_21_S_2_L_3_out, I0 =>  inp_feat(280), I1 =>  inp_feat(197), I2 =>  inp_feat(83), I3 =>  inp_feat(373), I4 =>  inp_feat(450), I5 =>  inp_feat(509)); 
C_21_S_2_L_4_inst : LUT6 generic map(INIT => "1000010101100101000101010001111110010011100100110001011111011111") port map( O =>C_21_S_2_L_4_out, I0 =>  inp_feat(65), I1 =>  inp_feat(210), I2 =>  inp_feat(83), I3 =>  inp_feat(449), I4 =>  inp_feat(185), I5 =>  inp_feat(35)); 
C_21_S_2_L_5_inst : LUT6 generic map(INIT => "0111111001000101011111000000111001010100011011000000111011001110") port map( O =>C_21_S_2_L_5_out, I0 =>  inp_feat(50), I1 =>  inp_feat(451), I2 =>  inp_feat(83), I3 =>  inp_feat(303), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_3_L_0_inst : LUT6 generic map(INIT => "1000000101001100000101000000110000100100111011000100110111001101") port map( O =>C_21_S_3_L_0_out, I0 =>  inp_feat(65), I1 =>  inp_feat(451), I2 =>  inp_feat(83), I3 =>  inp_feat(303), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_3_L_1_inst : LUT6 generic map(INIT => "0000110110011100001000101000110000100100010011000000110011101101") port map( O =>C_21_S_3_L_1_out, I0 =>  inp_feat(399), I1 =>  inp_feat(224), I2 =>  inp_feat(361), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_3_L_2_inst : LUT6 generic map(INIT => "1111111001111011100000110101011110010000110110110001011111111111") port map( O =>C_21_S_3_L_2_out, I0 =>  inp_feat(350), I1 =>  inp_feat(373), I2 =>  inp_feat(450), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_3_L_3_inst : LUT6 generic map(INIT => "0111110101001101100010100000000010011010000010001111100000000000") port map( O =>C_21_S_3_L_3_out, I0 =>  inp_feat(42), I1 =>  inp_feat(107), I2 =>  inp_feat(398), I3 =>  inp_feat(253), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_3_L_4_inst : LUT6 generic map(INIT => "0000010100010101000011010111111111000101100101110001011101111111") port map( O =>C_21_S_3_L_4_out, I0 =>  inp_feat(497), I1 =>  inp_feat(273), I2 =>  inp_feat(65), I3 =>  inp_feat(185), I4 =>  inp_feat(225), I5 =>  inp_feat(25)); 
C_21_S_3_L_5_inst : LUT6 generic map(INIT => "1011101110010111111000010001111110011001100111110001011111111111") port map( O =>C_21_S_3_L_5_out, I0 =>  inp_feat(210), I1 =>  inp_feat(65), I2 =>  inp_feat(450), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_4_L_0_inst : LUT6 generic map(INIT => "1010101110011100101000101000110000100100010011000000110011101101") port map( O =>C_21_S_4_L_0_out, I0 =>  inp_feat(399), I1 =>  inp_feat(224), I2 =>  inp_feat(361), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_4_L_1_inst : LUT6 generic map(INIT => "0100010000000010000000100010101110100110001101110010101011111111") port map( O =>C_21_S_4_L_1_out, I0 =>  inp_feat(15), I1 =>  inp_feat(112), I2 =>  inp_feat(361), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_4_L_2_inst : LUT6 generic map(INIT => "1010101110101011101000100010101001100000111010110010101110101011") port map( O =>C_21_S_4_L_2_out, I0 =>  inp_feat(346), I1 =>  inp_feat(65), I2 =>  inp_feat(450), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_4_L_3_inst : LUT6 generic map(INIT => "0100010110100110000000100010001010000000101010100010101010101010") port map( O =>C_21_S_4_L_3_out, I0 =>  inp_feat(253), I1 =>  inp_feat(350), I2 =>  inp_feat(83), I3 =>  inp_feat(303), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_4_L_4_inst : LUT6 generic map(INIT => "0110101011001110111001100100111001101100010011000100110011001100") port map( O =>C_21_S_4_L_4_out, I0 =>  inp_feat(215), I1 =>  inp_feat(230), I2 =>  inp_feat(65), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_4_L_5_inst : LUT6 generic map(INIT => "0110001000000000101010110000001011110011000001111011011100111011") port map( O =>C_21_S_4_L_5_out, I0 =>  inp_feat(358), I1 =>  inp_feat(454), I2 =>  inp_feat(384), I3 =>  inp_feat(227), I4 =>  inp_feat(175), I5 =>  inp_feat(405)); 
C_21_S_5_L_0_inst : LUT6 generic map(INIT => "1101110011011101011001100100110000000100010011100000000000001011") port map( O =>C_21_S_5_L_0_out, I0 =>  inp_feat(335), I1 =>  inp_feat(421), I2 =>  inp_feat(69), I3 =>  inp_feat(384), I4 =>  inp_feat(261), I5 =>  inp_feat(201)); 
C_21_S_5_L_1_inst : LUT6 generic map(INIT => "0000100100010100000000000000110000000000010011000000110011101101") port map( O =>C_21_S_5_L_1_out, I0 =>  inp_feat(399), I1 =>  inp_feat(224), I2 =>  inp_feat(361), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_5_L_2_inst : LUT6 generic map(INIT => "1000100000100100000011101011001110010000010000001010001011111010") port map( O =>C_21_S_5_L_2_out, I0 =>  inp_feat(435), I1 =>  inp_feat(26), I2 =>  inp_feat(66), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(388)); 
C_21_S_5_L_3_inst : LUT6 generic map(INIT => "0000000100100011001000100010101001100000011010110010101110101011") port map( O =>C_21_S_5_L_3_out, I0 =>  inp_feat(346), I1 =>  inp_feat(65), I2 =>  inp_feat(450), I3 =>  inp_feat(83), I4 =>  inp_feat(449), I5 =>  inp_feat(185)); 
C_21_S_5_L_4_inst : LUT6 generic map(INIT => "0000010010001000110110000000100001011100100010001110000010001000") port map( O =>C_21_S_5_L_4_out, I0 =>  inp_feat(84), I1 =>  inp_feat(189), I2 =>  inp_feat(361), I3 =>  inp_feat(185), I4 =>  inp_feat(130), I5 =>  inp_feat(422)); 
C_21_S_5_L_5_inst : LUT6 generic map(INIT => "1010100011000001111100000010000000111001010010000111100000111010") port map( O =>C_21_S_5_L_5_out, I0 =>  inp_feat(245), I1 =>  inp_feat(399), I2 =>  inp_feat(427), I3 =>  inp_feat(227), I4 =>  inp_feat(175), I5 =>  inp_feat(405)); 
C_22_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000111000000110011011100000001010111110001011111111111") port map( O =>C_22_S_0_L_0_out, I0 =>  inp_feat(83), I1 =>  inp_feat(350), I2 =>  inp_feat(399), I3 =>  inp_feat(324), I4 =>  inp_feat(373), I5 =>  inp_feat(185)); 
C_22_S_0_L_1_inst : LUT6 generic map(INIT => "0100000000000011111110110000101111111101000000001111110101000010") port map( O =>C_22_S_0_L_1_out, I0 =>  inp_feat(96), I1 =>  inp_feat(447), I2 =>  inp_feat(193), I3 =>  inp_feat(434), I4 =>  inp_feat(65), I5 =>  inp_feat(497)); 
C_22_S_0_L_2_inst : LUT6 generic map(INIT => "1110010100000011101101110010001110101110001000001011111010111010") port map( O =>C_22_S_0_L_2_out, I0 =>  inp_feat(278), I1 =>  inp_feat(160), I2 =>  inp_feat(468), I3 =>  inp_feat(119), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_22_S_0_L_3_inst : LUT6 generic map(INIT => "0000010011100000111100010000000011110001110100001111011100000000") port map( O =>C_22_S_0_L_3_out, I0 =>  inp_feat(83), I1 =>  inp_feat(61), I2 =>  inp_feat(316), I3 =>  inp_feat(253), I4 =>  inp_feat(280), I5 =>  inp_feat(112)); 
C_22_S_0_L_4_inst : LUT6 generic map(INIT => "1101111111111111000101000010110100000000100100000000000000000000") port map( O =>C_22_S_0_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(141), I2 =>  inp_feat(489), I3 =>  inp_feat(450), I4 =>  inp_feat(152), I5 =>  inp_feat(51)); 
C_22_S_0_L_5_inst : LUT6 generic map(INIT => "0000000100110011101110111101111110011101000111111001111111111111") port map( O =>C_22_S_0_L_5_out, I0 =>  inp_feat(497), I1 =>  inp_feat(288), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(361), I5 =>  inp_feat(35)); 
C_22_S_1_L_0_inst : LUT6 generic map(INIT => "0100000000000011111110110000101111111101000000001111110101000010") port map( O =>C_22_S_1_L_0_out, I0 =>  inp_feat(96), I1 =>  inp_feat(447), I2 =>  inp_feat(193), I3 =>  inp_feat(434), I4 =>  inp_feat(65), I5 =>  inp_feat(497)); 
C_22_S_1_L_1_inst : LUT6 generic map(INIT => "1110010100000011101101110010001110101110001000001011111010111010") port map( O =>C_22_S_1_L_1_out, I0 =>  inp_feat(278), I1 =>  inp_feat(160), I2 =>  inp_feat(468), I3 =>  inp_feat(119), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_22_S_1_L_2_inst : LUT6 generic map(INIT => "0000010011100000111100010000000011110001110100001111011100000000") port map( O =>C_22_S_1_L_2_out, I0 =>  inp_feat(83), I1 =>  inp_feat(61), I2 =>  inp_feat(316), I3 =>  inp_feat(253), I4 =>  inp_feat(280), I5 =>  inp_feat(112)); 
C_22_S_1_L_3_inst : LUT6 generic map(INIT => "1101111111111111000101000010110100000000100100000000000000000000") port map( O =>C_22_S_1_L_3_out, I0 =>  inp_feat(328), I1 =>  inp_feat(141), I2 =>  inp_feat(489), I3 =>  inp_feat(450), I4 =>  inp_feat(152), I5 =>  inp_feat(51)); 
C_22_S_1_L_4_inst : LUT6 generic map(INIT => "0000000100110011101110111101111110011101000111111001111111111111") port map( O =>C_22_S_1_L_4_out, I0 =>  inp_feat(497), I1 =>  inp_feat(288), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(361), I5 =>  inp_feat(35)); 
C_22_S_1_L_5_inst : LUT6 generic map(INIT => "1100100000000111001011111101111111000100001111111101111111111111") port map( O =>C_22_S_1_L_5_out, I0 =>  inp_feat(112), I1 =>  inp_feat(77), I2 =>  inp_feat(497), I3 =>  inp_feat(96), I4 =>  inp_feat(65), I5 =>  inp_feat(35)); 
C_22_S_2_L_0_inst : LUT6 generic map(INIT => "1000010001000100010011111111010001001100111101001100011111111100") port map( O =>C_22_S_2_L_0_out, I0 =>  inp_feat(65), I1 =>  inp_feat(66), I2 =>  inp_feat(468), I3 =>  inp_feat(280), I4 =>  inp_feat(328), I5 =>  inp_feat(35)); 
C_22_S_2_L_1_inst : LUT6 generic map(INIT => "0010000001111111010001111101111111001100110111110011111111111111") port map( O =>C_22_S_2_L_1_out, I0 =>  inp_feat(112), I1 =>  inp_feat(77), I2 =>  inp_feat(497), I3 =>  inp_feat(65), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_2_L_2_inst : LUT6 generic map(INIT => "1100100011000111000001111101111111000100110111110111111111111111") port map( O =>C_22_S_2_L_2_out, I0 =>  inp_feat(112), I1 =>  inp_feat(77), I2 =>  inp_feat(497), I3 =>  inp_feat(65), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_2_L_3_inst : LUT6 generic map(INIT => "0100000011010111011010001101111100011101110101110011111101111111") port map( O =>C_22_S_2_L_3_out, I0 =>  inp_feat(210), I1 =>  inp_feat(318), I2 =>  inp_feat(497), I3 =>  inp_feat(65), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_2_L_4_inst : LUT6 generic map(INIT => "1000111000101110111011100101110111100100011011010100110111111111") port map( O =>C_22_S_2_L_4_out, I0 =>  inp_feat(449), I1 =>  inp_feat(137), I2 =>  inp_feat(280), I3 =>  inp_feat(318), I4 =>  inp_feat(35), I5 =>  inp_feat(350)); 
C_22_S_2_L_5_inst : LUT6 generic map(INIT => "0110000000101110011010000110110010001000111011011100110111011101") port map( O =>C_22_S_2_L_5_out, I0 =>  inp_feat(185), I1 =>  inp_feat(456), I2 =>  inp_feat(305), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_3_L_0_inst : LUT6 generic map(INIT => "0111011001011111010001111101111101000100110111110011111111111111") port map( O =>C_22_S_3_L_0_out, I0 =>  inp_feat(112), I1 =>  inp_feat(77), I2 =>  inp_feat(497), I3 =>  inp_feat(65), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_3_L_1_inst : LUT6 generic map(INIT => "1010110100010100010111011111000101010100111101111111001111110111") port map( O =>C_22_S_3_L_1_out, I0 =>  inp_feat(361), I1 =>  inp_feat(497), I2 =>  inp_feat(468), I3 =>  inp_feat(318), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_22_S_3_L_2_inst : LUT6 generic map(INIT => "0000111101101111001100110111111111101001111111111001011101111111") port map( O =>C_22_S_3_L_2_out, I0 =>  inp_feat(83), I1 =>  inp_feat(303), I2 =>  inp_feat(210), I3 =>  inp_feat(65), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_3_L_3_inst : LUT6 generic map(INIT => "1101110000110101000111010011011111111101001111111101111111111111") port map( O =>C_22_S_3_L_3_out, I0 =>  inp_feat(65), I1 =>  inp_feat(83), I2 =>  inp_feat(318), I3 =>  inp_feat(280), I4 =>  inp_feat(35), I5 =>  inp_feat(350)); 
C_22_S_3_L_4_inst : LUT6 generic map(INIT => "0101000110011011001111110011111111010111110111110011011101111111") port map( O =>C_22_S_3_L_4_out, I0 =>  inp_feat(210), I1 =>  inp_feat(303), I2 =>  inp_feat(76), I3 =>  inp_feat(328), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_3_L_5_inst : LUT6 generic map(INIT => "0010100101110011011001001011000011111101000010000010001000100000") port map( O =>C_22_S_3_L_5_out, I0 =>  inp_feat(266), I1 =>  inp_feat(328), I2 =>  inp_feat(437), I3 =>  inp_feat(185), I4 =>  inp_feat(218), I5 =>  inp_feat(392)); 
C_22_S_4_L_0_inst : LUT6 generic map(INIT => "1011010110101001010011010110001111111111111100011111111100000101") port map( O =>C_22_S_4_L_0_out, I0 =>  inp_feat(361), I1 =>  inp_feat(93), I2 =>  inp_feat(26), I3 =>  inp_feat(456), I4 =>  inp_feat(303), I5 =>  inp_feat(280)); 
C_22_S_4_L_1_inst : LUT6 generic map(INIT => "0000001000101110111100101011001000111011001110101111000011110011") port map( O =>C_22_S_4_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(489), I2 =>  inp_feat(276), I3 =>  inp_feat(449), I4 =>  inp_feat(450), I5 =>  inp_feat(214)); 
C_22_S_4_L_2_inst : LUT6 generic map(INIT => "1101000101011111111101010111111111010101011111110011111111111111") port map( O =>C_22_S_4_L_2_out, I0 =>  inp_feat(65), I1 =>  inp_feat(91), I2 =>  inp_feat(305), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_4_L_3_inst : LUT6 generic map(INIT => "0111111111011110010000001100110011011010001011111000110011001101") port map( O =>C_22_S_4_L_3_out, I0 =>  inp_feat(95), I1 =>  inp_feat(307), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_4_L_4_inst : LUT6 generic map(INIT => "1110100110100010101011100010100000000100000000001100111101000000") port map( O =>C_22_S_4_L_4_out, I0 =>  inp_feat(110), I1 =>  inp_feat(128), I2 =>  inp_feat(141), I3 =>  inp_feat(144), I4 =>  inp_feat(29), I5 =>  inp_feat(304)); 
C_22_S_4_L_5_inst : LUT6 generic map(INIT => "0010000011010100001000100010000000000001000000100000000001000000") port map( O =>C_22_S_4_L_5_out, I0 =>  inp_feat(482), I1 =>  inp_feat(65), I2 =>  inp_feat(421), I3 =>  inp_feat(64), I4 =>  inp_feat(316), I5 =>  inp_feat(151)); 
C_22_S_5_L_0_inst : LUT6 generic map(INIT => "0000001011100110000001011101110110000110010111010000111011101111") port map( O =>C_22_S_5_L_0_out, I0 =>  inp_feat(289), I1 =>  inp_feat(137), I2 =>  inp_feat(318), I3 =>  inp_feat(280), I4 =>  inp_feat(35), I5 =>  inp_feat(350)); 
C_22_S_5_L_1_inst : LUT6 generic map(INIT => "1111110111010111001010011111111100110111111101110011011111111111") port map( O =>C_22_S_5_L_1_out, I0 =>  inp_feat(272), I1 =>  inp_feat(318), I2 =>  inp_feat(76), I3 =>  inp_feat(303), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_5_L_2_inst : LUT6 generic map(INIT => "0000100100101000110001001000100010001110000110101000100010001010") port map( O =>C_22_S_5_L_2_out, I0 =>  inp_feat(94), I1 =>  inp_feat(307), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_22_S_5_L_3_inst : LUT6 generic map(INIT => "0111011111000011000101110000100111100111101000001110011110000001") port map( O =>C_22_S_5_L_3_out, I0 =>  inp_feat(450), I1 =>  inp_feat(497), I2 =>  inp_feat(280), I3 =>  inp_feat(182), I4 =>  inp_feat(25), I5 =>  inp_feat(29)); 
C_22_S_5_L_4_inst : LUT6 generic map(INIT => "1101100111011101000000011100000011111101111101110001000011000000") port map( O =>C_22_S_5_L_4_out, I0 =>  inp_feat(201), I1 =>  inp_feat(281), I2 =>  inp_feat(142), I3 =>  inp_feat(392), I4 =>  inp_feat(425), I5 =>  inp_feat(391)); 
C_22_S_5_L_5_inst : LUT6 generic map(INIT => "0011001010110010000000001101000111001101101000000000101011000000") port map( O =>C_22_S_5_L_5_out, I0 =>  inp_feat(81), I1 =>  inp_feat(64), I2 =>  inp_feat(57), I3 =>  inp_feat(188), I4 =>  inp_feat(435), I5 =>  inp_feat(391)); 
C_23_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000111000000010101011100000001001101110001011101111111") port map( O =>C_23_S_0_L_0_out, I0 =>  inp_feat(350), I1 =>  inp_feat(83), I2 =>  inp_feat(399), I3 =>  inp_feat(324), I4 =>  inp_feat(373), I5 =>  inp_feat(185)); 
C_23_S_0_L_1_inst : LUT6 generic map(INIT => "0010000100111000001101011111000010111000101100001111000011110001") port map( O =>C_23_S_0_L_1_out, I0 =>  inp_feat(112), I1 =>  inp_feat(35), I2 =>  inp_feat(245), I3 =>  inp_feat(210), I4 =>  inp_feat(65), I5 =>  inp_feat(497)); 
C_23_S_0_L_2_inst : LUT6 generic map(INIT => "1101000110111110111100010000000000000000000110101000000000010000") port map( O =>C_23_S_0_L_2_out, I0 =>  inp_feat(296), I1 =>  inp_feat(509), I2 =>  inp_feat(280), I3 =>  inp_feat(318), I4 =>  inp_feat(11), I5 =>  inp_feat(183)); 
C_23_S_0_L_3_inst : LUT6 generic map(INIT => "0000001000000100110000011010101100100010000010111100100010000000") port map( O =>C_23_S_0_L_3_out, I0 =>  inp_feat(321), I1 =>  inp_feat(385), I2 =>  inp_feat(463), I3 =>  inp_feat(245), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_0_L_4_inst : LUT6 generic map(INIT => "1110011100000101011011100000000011111111101011111100111100001110") port map( O =>C_23_S_0_L_4_out, I0 =>  inp_feat(431), I1 =>  inp_feat(126), I2 =>  inp_feat(471), I3 =>  inp_feat(251), I4 =>  inp_feat(29), I5 =>  inp_feat(283)); 
C_23_S_0_L_5_inst : LUT6 generic map(INIT => "1000100000010000101000010000000000111000000010001011001000000000") port map( O =>C_23_S_0_L_5_out, I0 =>  inp_feat(138), I1 =>  inp_feat(449), I2 =>  inp_feat(463), I3 =>  inp_feat(245), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_1_L_0_inst : LUT6 generic map(INIT => "0010000100111000001101011111000010111000101100001111000011110001") port map( O =>C_23_S_1_L_0_out, I0 =>  inp_feat(112), I1 =>  inp_feat(35), I2 =>  inp_feat(245), I3 =>  inp_feat(210), I4 =>  inp_feat(65), I5 =>  inp_feat(497)); 
C_23_S_1_L_1_inst : LUT6 generic map(INIT => "1101000110111110111100010000000000000000000110101000000000010000") port map( O =>C_23_S_1_L_1_out, I0 =>  inp_feat(296), I1 =>  inp_feat(509), I2 =>  inp_feat(280), I3 =>  inp_feat(318), I4 =>  inp_feat(11), I5 =>  inp_feat(183)); 
C_23_S_1_L_2_inst : LUT6 generic map(INIT => "0000001000000100110000011010101100100010000010111100100010000000") port map( O =>C_23_S_1_L_2_out, I0 =>  inp_feat(321), I1 =>  inp_feat(385), I2 =>  inp_feat(463), I3 =>  inp_feat(245), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_1_L_3_inst : LUT6 generic map(INIT => "1110011100000101011011100000000011111111101011111100111100001110") port map( O =>C_23_S_1_L_3_out, I0 =>  inp_feat(431), I1 =>  inp_feat(126), I2 =>  inp_feat(471), I3 =>  inp_feat(251), I4 =>  inp_feat(29), I5 =>  inp_feat(283)); 
C_23_S_1_L_4_inst : LUT6 generic map(INIT => "1000100000010000101000010000000000111000000010001011001000000000") port map( O =>C_23_S_1_L_4_out, I0 =>  inp_feat(138), I1 =>  inp_feat(449), I2 =>  inp_feat(463), I3 =>  inp_feat(245), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_1_L_5_inst : LUT6 generic map(INIT => "0001000100010001000010001000000001011100011000101000101000000000") port map( O =>C_23_S_1_L_5_out, I0 =>  inp_feat(334), I1 =>  inp_feat(180), I2 =>  inp_feat(210), I3 =>  inp_feat(307), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_2_L_0_inst : LUT6 generic map(INIT => "1111100110001100111100000100000000000001000011000011000100010000") port map( O =>C_23_S_2_L_0_out, I0 =>  inp_feat(316), I1 =>  inp_feat(317), I2 =>  inp_feat(65), I3 =>  inp_feat(83), I4 =>  inp_feat(11), I5 =>  inp_feat(183)); 
C_23_S_2_L_1_inst : LUT6 generic map(INIT => "1000111110000000000000001000100001110010100010001000000010101000") port map( O =>C_23_S_2_L_1_out, I0 =>  inp_feat(413), I1 =>  inp_feat(248), I2 =>  inp_feat(403), I3 =>  inp_feat(318), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_2_L_2_inst : LUT6 generic map(INIT => "0001010100000000100000010000010010010010000001101100110000000000") port map( O =>C_23_S_2_L_2_out, I0 =>  inp_feat(468), I1 =>  inp_feat(385), I2 =>  inp_feat(463), I3 =>  inp_feat(245), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_2_L_3_inst : LUT6 generic map(INIT => "1100010010100000011110010000000011111011101110111111110001010101") port map( O =>C_23_S_2_L_3_out, I0 =>  inp_feat(464), I1 =>  inp_feat(321), I2 =>  inp_feat(486), I3 =>  inp_feat(101), I4 =>  inp_feat(29), I5 =>  inp_feat(283)); 
C_23_S_2_L_4_inst : LUT6 generic map(INIT => "0000011111011111000101110111111111001000000000000000000000000000") port map( O =>C_23_S_2_L_4_out, I0 =>  inp_feat(272), I1 =>  inp_feat(450), I2 =>  inp_feat(318), I3 =>  inp_feat(280), I4 =>  inp_feat(35), I5 =>  inp_feat(283)); 
C_23_S_2_L_5_inst : LUT6 generic map(INIT => "1001010100101100001100111000000001010111111000001111111100000000") port map( O =>C_23_S_2_L_5_out, I0 =>  inp_feat(318), I1 =>  inp_feat(35), I2 =>  inp_feat(115), I3 =>  inp_feat(81), I4 =>  inp_feat(497), I5 =>  inp_feat(65)); 
C_23_S_3_L_0_inst : LUT6 generic map(INIT => "1110001001100100000001000110110000110110111111000100110011001100") port map( O =>C_23_S_3_L_0_out, I0 =>  inp_feat(318), I1 =>  inp_feat(317), I2 =>  inp_feat(83), I3 =>  inp_feat(65), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_3_L_1_inst : LUT6 generic map(INIT => "0000000011110100010001000110110010010110111111000100110001001100") port map( O =>C_23_S_3_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(317), I2 =>  inp_feat(83), I3 =>  inp_feat(65), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_3_L_2_inst : LUT6 generic map(INIT => "0000100110101000001000001010001011111101100001000101011000000000") port map( O =>C_23_S_3_L_2_out, I0 =>  inp_feat(334), I1 =>  inp_feat(210), I2 =>  inp_feat(180), I3 =>  inp_feat(318), I4 =>  inp_feat(35), I5 =>  inp_feat(277)); 
C_23_S_3_L_3_inst : LUT6 generic map(INIT => "1100010000010011000111101001111101010011101101110111111101111111") port map( O =>C_23_S_3_L_3_out, I0 =>  inp_feat(93), I1 =>  inp_feat(318), I2 =>  inp_feat(13), I3 =>  inp_feat(160), I4 =>  inp_feat(303), I5 =>  inp_feat(280)); 
C_23_S_3_L_4_inst : LUT6 generic map(INIT => "0000100000111001011100100001101010101000000000001010000000000000") port map( O =>C_23_S_3_L_4_out, I0 =>  inp_feat(104), I1 =>  inp_feat(441), I2 =>  inp_feat(205), I3 =>  inp_feat(417), I4 =>  inp_feat(303), I5 =>  inp_feat(280)); 
C_23_S_3_L_5_inst : LUT6 generic map(INIT => "1111101111011110001010101110000000001111010101000000001100100000") port map( O =>C_23_S_3_L_5_out, I0 =>  inp_feat(190), I1 =>  inp_feat(72), I2 =>  inp_feat(132), I3 =>  inp_feat(456), I4 =>  inp_feat(251), I5 =>  inp_feat(29)); 
C_23_S_4_L_0_inst : LUT6 generic map(INIT => "0000000011010000000100001111000110100000110100011111000011110001") port map( O =>C_23_S_4_L_0_out, I0 =>  inp_feat(450), I1 =>  inp_feat(361), I2 =>  inp_feat(180), I3 =>  inp_feat(280), I4 =>  inp_feat(26), I5 =>  inp_feat(404)); 
C_23_S_4_L_1_inst : LUT6 generic map(INIT => "1010110000011011001000010000100100111000000010001011001000000000") port map( O =>C_23_S_4_L_1_out, I0 =>  inp_feat(138), I1 =>  inp_feat(449), I2 =>  inp_feat(463), I3 =>  inp_feat(245), I4 =>  inp_feat(280), I5 =>  inp_feat(35)); 
C_23_S_4_L_2_inst : LUT6 generic map(INIT => "0010010000100111000000010011011111001101001111110011011111111111") port map( O =>C_23_S_4_L_2_out, I0 =>  inp_feat(65), I1 =>  inp_feat(324), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_23_S_4_L_3_inst : LUT6 generic map(INIT => "1111110011011010111101001001100000000000110000101011000110101000") port map( O =>C_23_S_4_L_3_out, I0 =>  inp_feat(494), I1 =>  inp_feat(292), I2 =>  inp_feat(242), I3 =>  inp_feat(460), I4 =>  inp_feat(231), I5 =>  inp_feat(405)); 
C_23_S_4_L_4_inst : LUT6 generic map(INIT => "0100000000000111000000000011111100001101010111110011010101111111") port map( O =>C_23_S_4_L_4_out, I0 =>  inp_feat(361), I1 =>  inp_feat(324), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_23_S_4_L_5_inst : LUT6 generic map(INIT => "1001000111000010000111110000001010001011000000001001111100001101") port map( O =>C_23_S_4_L_5_out, I0 =>  inp_feat(160), I1 =>  inp_feat(56), I2 =>  inp_feat(462), I3 =>  inp_feat(96), I4 =>  inp_feat(261), I5 =>  inp_feat(47)); 
C_23_S_5_L_0_inst : LUT6 generic map(INIT => "0001100100011000011101010011100011000001100010000000000111100000") port map( O =>C_23_S_5_L_0_out, I0 =>  inp_feat(361), I1 =>  inp_feat(225), I2 =>  inp_feat(121), I3 =>  inp_feat(471), I4 =>  inp_feat(101), I5 =>  inp_feat(467)); 
C_23_S_5_L_1_inst : LUT6 generic map(INIT => "1001011111010111100010110000011101000001000001110100010100000011") port map( O =>C_23_S_5_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(83), I2 =>  inp_feat(361), I3 =>  inp_feat(29), I4 =>  inp_feat(486), I5 =>  inp_feat(467)); 
C_23_S_5_L_2_inst : LUT6 generic map(INIT => "1000100100010011100100010111111100010111010111110101111111111111") port map( O =>C_23_S_5_L_2_out, I0 =>  inp_feat(303), I1 =>  inp_feat(288), I2 =>  inp_feat(318), I3 =>  inp_feat(210), I4 =>  inp_feat(65), I5 =>  inp_feat(35)); 
C_23_S_5_L_3_inst : LUT6 generic map(INIT => "0000001001101011000000000010101100001000001011110010101010111111") port map( O =>C_23_S_5_L_3_out, I0 =>  inp_feat(183), I1 =>  inp_feat(324), I2 =>  inp_feat(210), I3 =>  inp_feat(318), I4 =>  inp_feat(96), I5 =>  inp_feat(35)); 
C_23_S_5_L_4_inst : LUT6 generic map(INIT => "1000100011100000100000100010000011101110001011000111111101000110") port map( O =>C_23_S_5_L_4_out, I0 =>  inp_feat(319), I1 =>  inp_feat(310), I2 =>  inp_feat(169), I3 =>  inp_feat(350), I4 =>  inp_feat(275), I5 =>  inp_feat(10)); 
C_23_S_5_L_5_inst : LUT6 generic map(INIT => "1000000101000111000111110111111111111001000000010000010100000111") port map( O =>C_23_S_5_L_5_out, I0 =>  inp_feat(210), I1 =>  inp_feat(449), I2 =>  inp_feat(83), I3 =>  inp_feat(221), I4 =>  inp_feat(445), I5 =>  inp_feat(130)); 
C_24_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111101010100011111111111000001111100010000000") port map( O =>C_24_S_0_L_0_out, I0 =>  inp_feat(18), I1 =>  inp_feat(67), I2 =>  inp_feat(389), I3 =>  inp_feat(421), I4 =>  inp_feat(354), I5 =>  inp_feat(287)); 
C_24_S_0_L_1_inst : LUT6 generic map(INIT => "1111111111101111010111110000110100000001001011110001111000001101") port map( O =>C_24_S_0_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(188), I2 =>  inp_feat(179), I3 =>  inp_feat(123), I4 =>  inp_feat(445), I5 =>  inp_feat(127)); 
C_24_S_0_L_2_inst : LUT6 generic map(INIT => "1110111000011010111100000010001011110010010110100010001001100010") port map( O =>C_24_S_0_L_2_out, I0 =>  inp_feat(174), I1 =>  inp_feat(31), I2 =>  inp_feat(195), I3 =>  inp_feat(423), I4 =>  inp_feat(94), I5 =>  inp_feat(169)); 
C_24_S_0_L_3_inst : LUT6 generic map(INIT => "1001011100010011110111111111001111111111111111001110110000001101") port map( O =>C_24_S_0_L_3_out, I0 =>  inp_feat(81), I1 =>  inp_feat(287), I2 =>  inp_feat(445), I3 =>  inp_feat(309), I4 =>  inp_feat(355), I5 =>  inp_feat(15)); 
C_24_S_0_L_4_inst : LUT6 generic map(INIT => "0010101001111110111111010110111000100110001000101111111111101010") port map( O =>C_24_S_0_L_4_out, I0 =>  inp_feat(67), I1 =>  inp_feat(331), I2 =>  inp_feat(120), I3 =>  inp_feat(244), I4 =>  inp_feat(170), I5 =>  inp_feat(72)); 
C_24_S_0_L_5_inst : LUT6 generic map(INIT => "1111010111011101111011101111111101000111111111111111001111111001") port map( O =>C_24_S_0_L_5_out, I0 =>  inp_feat(405), I1 =>  inp_feat(204), I2 =>  inp_feat(42), I3 =>  inp_feat(0), I4 =>  inp_feat(445), I5 =>  inp_feat(72)); 
C_24_S_1_L_0_inst : LUT6 generic map(INIT => "1111111111101111010111110000110100000001001011110001111000001101") port map( O =>C_24_S_1_L_0_out, I0 =>  inp_feat(44), I1 =>  inp_feat(188), I2 =>  inp_feat(179), I3 =>  inp_feat(123), I4 =>  inp_feat(445), I5 =>  inp_feat(127)); 
C_24_S_1_L_1_inst : LUT6 generic map(INIT => "1110111000011010111100000010001011110010010110100010001001100010") port map( O =>C_24_S_1_L_1_out, I0 =>  inp_feat(174), I1 =>  inp_feat(31), I2 =>  inp_feat(195), I3 =>  inp_feat(423), I4 =>  inp_feat(94), I5 =>  inp_feat(169)); 
C_24_S_1_L_2_inst : LUT6 generic map(INIT => "1001011100010011110111111111001111111111111111001110110000001101") port map( O =>C_24_S_1_L_2_out, I0 =>  inp_feat(81), I1 =>  inp_feat(287), I2 =>  inp_feat(445), I3 =>  inp_feat(309), I4 =>  inp_feat(355), I5 =>  inp_feat(15)); 
C_24_S_1_L_3_inst : LUT6 generic map(INIT => "0010101001111110111111010110111000100110001000101111111111101010") port map( O =>C_24_S_1_L_3_out, I0 =>  inp_feat(67), I1 =>  inp_feat(331), I2 =>  inp_feat(120), I3 =>  inp_feat(244), I4 =>  inp_feat(170), I5 =>  inp_feat(72)); 
C_24_S_1_L_4_inst : LUT6 generic map(INIT => "1111010111011101111011101111111101000111111111111111001111111001") port map( O =>C_24_S_1_L_4_out, I0 =>  inp_feat(405), I1 =>  inp_feat(204), I2 =>  inp_feat(42), I3 =>  inp_feat(0), I4 =>  inp_feat(445), I5 =>  inp_feat(72)); 
C_24_S_1_L_5_inst : LUT6 generic map(INIT => "1001010110011100111101111011010001010100110110001111110110000000") port map( O =>C_24_S_1_L_5_out, I0 =>  inp_feat(241), I1 =>  inp_feat(354), I2 =>  inp_feat(167), I3 =>  inp_feat(3), I4 =>  inp_feat(507), I5 =>  inp_feat(135)); 
C_24_S_2_L_0_inst : LUT6 generic map(INIT => "1011111111111111101010111010111000000101011101010010001100001010") port map( O =>C_24_S_2_L_0_out, I0 =>  inp_feat(46), I1 =>  inp_feat(279), I2 =>  inp_feat(371), I3 =>  inp_feat(284), I4 =>  inp_feat(127), I5 =>  inp_feat(169)); 
C_24_S_2_L_1_inst : LUT6 generic map(INIT => "0100000111111100011100011111011011101110111111111111010011111111") port map( O =>C_24_S_2_L_1_out, I0 =>  inp_feat(207), I1 =>  inp_feat(90), I2 =>  inp_feat(124), I3 =>  inp_feat(437), I4 =>  inp_feat(232), I5 =>  inp_feat(52)); 
C_24_S_2_L_2_inst : LUT6 generic map(INIT => "1101100001101110010111001110011011111010111011101111100001001000") port map( O =>C_24_S_2_L_2_out, I0 =>  inp_feat(287), I1 =>  inp_feat(94), I2 =>  inp_feat(169), I3 =>  inp_feat(115), I4 =>  inp_feat(75), I5 =>  inp_feat(12)); 
C_24_S_2_L_3_inst : LUT6 generic map(INIT => "1111101111111110111110101111110111111011011011110000000100111110") port map( O =>C_24_S_2_L_3_out, I0 =>  inp_feat(27), I1 =>  inp_feat(313), I2 =>  inp_feat(90), I3 =>  inp_feat(284), I4 =>  inp_feat(510), I5 =>  inp_feat(423)); 
C_24_S_2_L_4_inst : LUT6 generic map(INIT => "1110100100100011001000001110101101010011111110110000000010110000") port map( O =>C_24_S_2_L_4_out, I0 =>  inp_feat(427), I1 =>  inp_feat(172), I2 =>  inp_feat(275), I3 =>  inp_feat(371), I4 =>  inp_feat(20), I5 =>  inp_feat(187)); 
C_24_S_2_L_5_inst : LUT6 generic map(INIT => "0110001011000000111011101110100000000101000010001110111011000000") port map( O =>C_24_S_2_L_5_out, I0 =>  inp_feat(287), I1 =>  inp_feat(37), I2 =>  inp_feat(440), I3 =>  inp_feat(475), I4 =>  inp_feat(12), I5 =>  inp_feat(25)); 
C_24_S_3_L_0_inst : LUT6 generic map(INIT => "0000000011100110110101110110111011101110111011101010001011101000") port map( O =>C_24_S_3_L_0_out, I0 =>  inp_feat(287), I1 =>  inp_feat(261), I2 =>  inp_feat(394), I3 =>  inp_feat(437), I4 =>  inp_feat(232), I5 =>  inp_feat(52)); 
C_24_S_3_L_1_inst : LUT6 generic map(INIT => "1101011101111111101000011111111011010001111101100001001111111101") port map( O =>C_24_S_3_L_1_out, I0 =>  inp_feat(204), I1 =>  inp_feat(343), I2 =>  inp_feat(422), I3 =>  inp_feat(139), I4 =>  inp_feat(429), I5 =>  inp_feat(25)); 
C_24_S_3_L_2_inst : LUT6 generic map(INIT => "1111100110101101110010011101110010111100010010100101000011010000") port map( O =>C_24_S_3_L_2_out, I0 =>  inp_feat(321), I1 =>  inp_feat(503), I2 =>  inp_feat(94), I3 =>  inp_feat(81), I4 =>  inp_feat(287), I5 =>  inp_feat(140)); 
C_24_S_3_L_3_inst : LUT6 generic map(INIT => "1011100100101011101000100111111101001010000011001100111110001110") port map( O =>C_24_S_3_L_3_out, I0 =>  inp_feat(72), I1 =>  inp_feat(67), I2 =>  inp_feat(91), I3 =>  inp_feat(354), I4 =>  inp_feat(263), I5 =>  inp_feat(261)); 
C_24_S_3_L_4_inst : LUT6 generic map(INIT => "0000000000100110001100111111000111101110111011101111101110011011") port map( O =>C_24_S_3_L_4_out, I0 =>  inp_feat(127), I1 =>  inp_feat(20), I2 =>  inp_feat(510), I3 =>  inp_feat(44), I4 =>  inp_feat(1), I5 =>  inp_feat(241)); 
C_24_S_3_L_5_inst : LUT6 generic map(INIT => "1111100111110001101111101100010000010101111101101111111100101100") port map( O =>C_24_S_3_L_5_out, I0 =>  inp_feat(407), I1 =>  inp_feat(4), I2 =>  inp_feat(320), I3 =>  inp_feat(338), I4 =>  inp_feat(5), I5 =>  inp_feat(151)); 
C_24_S_4_L_0_inst : LUT6 generic map(INIT => "0010101010001110010111101111111011011111111111010110100011110000") port map( O =>C_24_S_4_L_0_out, I0 =>  inp_feat(180), I1 =>  inp_feat(27), I2 =>  inp_feat(23), I3 =>  inp_feat(347), I4 =>  inp_feat(129), I5 =>  inp_feat(391)); 
C_24_S_4_L_1_inst : LUT6 generic map(INIT => "1111101010111000101101111110101000111111101100001111101110101010") port map( O =>C_24_S_4_L_1_out, I0 =>  inp_feat(501), I1 =>  inp_feat(478), I2 =>  inp_feat(99), I3 =>  inp_feat(342), I4 =>  inp_feat(263), I5 =>  inp_feat(261)); 
C_24_S_4_L_2_inst : LUT6 generic map(INIT => "0000011000011100011011100101100011101100111111101010000000101000") port map( O =>C_24_S_4_L_2_out, I0 =>  inp_feat(287), I1 =>  inp_feat(67), I2 =>  inp_feat(501), I3 =>  inp_feat(325), I4 =>  inp_feat(320), I5 =>  inp_feat(74)); 
C_24_S_4_L_3_inst : LUT6 generic map(INIT => "1101100111011100001111011100110000010000110111000011010011000100") port map( O =>C_24_S_4_L_3_out, I0 =>  inp_feat(91), I1 =>  inp_feat(354), I2 =>  inp_feat(475), I3 =>  inp_feat(68), I4 =>  inp_feat(125), I5 =>  inp_feat(25)); 
C_24_S_4_L_4_inst : LUT6 generic map(INIT => "0110101010101000011000101111100011111110111100001111110000000000") port map( O =>C_24_S_4_L_4_out, I0 =>  inp_feat(46), I1 =>  inp_feat(354), I2 =>  inp_feat(94), I3 =>  inp_feat(50), I4 =>  inp_feat(44), I5 =>  inp_feat(291)); 
C_24_S_4_L_5_inst : LUT6 generic map(INIT => "1101001100100111101111111111011011000100110111001100110011001000") port map( O =>C_24_S_4_L_5_out, I0 =>  inp_feat(453), I1 =>  inp_feat(45), I2 =>  inp_feat(429), I3 =>  inp_feat(232), I4 =>  inp_feat(288), I5 =>  inp_feat(220)); 
C_24_S_5_L_0_inst : LUT6 generic map(INIT => "0100011110100100000111001101110011111000111111111111111111111111") port map( O =>C_24_S_5_L_0_out, I0 =>  inp_feat(92), I1 =>  inp_feat(277), I2 =>  inp_feat(426), I3 =>  inp_feat(232), I4 =>  inp_feat(288), I5 =>  inp_feat(220)); 
C_24_S_5_L_1_inst : LUT6 generic map(INIT => "1110110011101000000011101110100000101110111111110000100010100000") port map( O =>C_24_S_5_L_1_out, I0 =>  inp_feat(152), I1 =>  inp_feat(155), I2 =>  inp_feat(420), I3 =>  inp_feat(1), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_24_S_5_L_2_inst : LUT6 generic map(INIT => "1010101011100110011101101110100011001100010011000001010011000000") port map( O =>C_24_S_5_L_2_out, I0 =>  inp_feat(287), I1 =>  inp_feat(67), I2 =>  inp_feat(261), I3 =>  inp_feat(158), I4 =>  inp_feat(403), I5 =>  inp_feat(113)); 
C_24_S_5_L_3_inst : LUT6 generic map(INIT => "1001010111110111111111011111011100010001100000101111111100110111") port map( O =>C_24_S_5_L_3_out, I0 =>  inp_feat(256), I1 =>  inp_feat(395), I2 =>  inp_feat(415), I3 =>  inp_feat(313), I4 =>  inp_feat(172), I5 =>  inp_feat(100)); 
C_24_S_5_L_4_inst : LUT6 generic map(INIT => "0011101101101011011011111010101111111110011111111111111110101011") port map( O =>C_24_S_5_L_4_out, I0 =>  inp_feat(321), I1 =>  inp_feat(339), I2 =>  inp_feat(327), I3 =>  inp_feat(389), I4 =>  inp_feat(71), I5 =>  inp_feat(203)); 
C_24_S_5_L_5_inst : LUT6 generic map(INIT => "1111110111111110111100101111110101011011101111101111010110101011") port map( O =>C_24_S_5_L_5_out, I0 =>  inp_feat(139), I1 =>  inp_feat(378), I2 =>  inp_feat(321), I3 =>  inp_feat(87), I4 =>  inp_feat(105), I5 =>  inp_feat(43)); 
C_25_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000000000000000000011100000000000101110001001101111111") port map( O =>C_25_S_0_L_0_out, I0 =>  inp_feat(127), I1 =>  inp_feat(67), I2 =>  inp_feat(389), I3 =>  inp_feat(421), I4 =>  inp_feat(354), I5 =>  inp_feat(287)); 
C_25_S_0_L_1_inst : LUT6 generic map(INIT => "0000000011100100101110111110000111111000101000001110000011110000") port map( O =>C_25_S_0_L_1_out, I0 =>  inp_feat(90), I1 =>  inp_feat(81), I2 =>  inp_feat(342), I3 =>  inp_feat(127), I4 =>  inp_feat(46), I5 =>  inp_feat(121)); 
C_25_S_0_L_2_inst : LUT6 generic map(INIT => "1110110010000000100010000000000000001010000000110000010000000000") port map( O =>C_25_S_0_L_2_out, I0 =>  inp_feat(375), I1 =>  inp_feat(81), I2 =>  inp_feat(9), I3 =>  inp_feat(312), I4 =>  inp_feat(32), I5 =>  inp_feat(98)); 
C_25_S_0_L_3_inst : LUT6 generic map(INIT => "0100010000010001000001001100000011101110100001010100000000000010") port map( O =>C_25_S_0_L_3_out, I0 =>  inp_feat(195), I1 =>  inp_feat(317), I2 =>  inp_feat(2), I3 =>  inp_feat(151), I4 =>  inp_feat(397), I5 =>  inp_feat(303)); 
C_25_S_0_L_4_inst : LUT6 generic map(INIT => "1110001010100010110111110000000011110110000010001111111100000100") port map( O =>C_25_S_0_L_4_out, I0 =>  inp_feat(287), I1 =>  inp_feat(44), I2 =>  inp_feat(67), I3 =>  inp_feat(17), I4 =>  inp_feat(421), I5 =>  inp_feat(107)); 
C_25_S_0_L_5_inst : LUT6 generic map(INIT => "0001000111010000010100010100000110111011100000000111111100000001") port map( O =>C_25_S_0_L_5_out, I0 =>  inp_feat(67), I1 =>  inp_feat(94), I2 =>  inp_feat(46), I3 =>  inp_feat(279), I4 =>  inp_feat(261), I5 =>  inp_feat(354)); 
C_25_S_1_L_0_inst : LUT6 generic map(INIT => "0000000011100100101110111110000111111000101000001110000011110000") port map( O =>C_25_S_1_L_0_out, I0 =>  inp_feat(90), I1 =>  inp_feat(81), I2 =>  inp_feat(342), I3 =>  inp_feat(127), I4 =>  inp_feat(46), I5 =>  inp_feat(121)); 
C_25_S_1_L_1_inst : LUT6 generic map(INIT => "1110110010000000100010000000000000001010000000110000010000000000") port map( O =>C_25_S_1_L_1_out, I0 =>  inp_feat(375), I1 =>  inp_feat(81), I2 =>  inp_feat(9), I3 =>  inp_feat(312), I4 =>  inp_feat(32), I5 =>  inp_feat(98)); 
C_25_S_1_L_2_inst : LUT6 generic map(INIT => "0100010000010001000001001100000011101110100001010100000000000010") port map( O =>C_25_S_1_L_2_out, I0 =>  inp_feat(195), I1 =>  inp_feat(317), I2 =>  inp_feat(2), I3 =>  inp_feat(151), I4 =>  inp_feat(397), I5 =>  inp_feat(303)); 
C_25_S_1_L_3_inst : LUT6 generic map(INIT => "1110001010100010110111110000000011110110000010001111111100000100") port map( O =>C_25_S_1_L_3_out, I0 =>  inp_feat(287), I1 =>  inp_feat(44), I2 =>  inp_feat(67), I3 =>  inp_feat(17), I4 =>  inp_feat(421), I5 =>  inp_feat(107)); 
C_25_S_1_L_4_inst : LUT6 generic map(INIT => "0001000111010000010100010100000110111011100000000111111100000001") port map( O =>C_25_S_1_L_4_out, I0 =>  inp_feat(67), I1 =>  inp_feat(94), I2 =>  inp_feat(46), I3 =>  inp_feat(279), I4 =>  inp_feat(261), I5 =>  inp_feat(354)); 
C_25_S_1_L_5_inst : LUT6 generic map(INIT => "1011011100000000111101101110010000100000000000001110100011100000") port map( O =>C_25_S_1_L_5_out, I0 =>  inp_feat(491), I1 =>  inp_feat(288), I2 =>  inp_feat(106), I3 =>  inp_feat(277), I4 =>  inp_feat(0), I5 =>  inp_feat(256)); 
C_25_S_2_L_0_inst : LUT6 generic map(INIT => "1010010000101011100100010111111110110110111111110011110101111111") port map( O =>C_25_S_2_L_0_out, I0 =>  inp_feat(287), I1 =>  inp_feat(304), I2 =>  inp_feat(428), I3 =>  inp_feat(354), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_25_S_2_L_1_inst : LUT6 generic map(INIT => "0001000010001001111000000001000010111011100100000111011110010000") port map( O =>C_25_S_2_L_1_out, I0 =>  inp_feat(421), I1 =>  inp_feat(94), I2 =>  inp_feat(476), I3 =>  inp_feat(277), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_2_L_2_inst : LUT6 generic map(INIT => "1000000001101100001001000100110010010110011011000110110011001101") port map( O =>C_25_S_2_L_2_out, I0 =>  inp_feat(94), I1 =>  inp_feat(279), I2 =>  inp_feat(503), I3 =>  inp_feat(354), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_25_S_2_L_3_inst : LUT6 generic map(INIT => "1001000011100000111010001110001100000000100000001011000000000000") port map( O =>C_25_S_2_L_3_out, I0 =>  inp_feat(221), I1 =>  inp_feat(397), I2 =>  inp_feat(145), I3 =>  inp_feat(306), I4 =>  inp_feat(325), I5 =>  inp_feat(57)); 
C_25_S_2_L_4_inst : LUT6 generic map(INIT => "0000001000000000100011010010001001000000111100001010000010110010") port map( O =>C_25_S_2_L_4_out, I0 =>  inp_feat(262), I1 =>  inp_feat(94), I2 =>  inp_feat(385), I3 =>  inp_feat(46), I4 =>  inp_feat(261), I5 =>  inp_feat(354)); 
C_25_S_2_L_5_inst : LUT6 generic map(INIT => "1010101101110100110111011100100100000000000100011100100010000000") port map( O =>C_25_S_2_L_5_out, I0 =>  inp_feat(106), I1 =>  inp_feat(499), I2 =>  inp_feat(73), I3 =>  inp_feat(48), I4 =>  inp_feat(112), I5 =>  inp_feat(99)); 
C_25_S_3_L_0_inst : LUT6 generic map(INIT => "1000010100001111000100010001011100000011101111110111111101011111") port map( O =>C_25_S_3_L_0_out, I0 =>  inp_feat(354), I1 =>  inp_feat(18), I2 =>  inp_feat(503), I3 =>  inp_feat(183), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_3_L_1_inst : LUT6 generic map(INIT => "0001001001010011100000011010001101001010011111110001011101111111") port map( O =>C_25_S_3_L_1_out, I0 =>  inp_feat(127), I1 =>  inp_feat(67), I2 =>  inp_feat(94), I3 =>  inp_feat(140), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_3_L_2_inst : LUT6 generic map(INIT => "1011110010100001100100000000000011011100000000001110110111000000") port map( O =>C_25_S_3_L_2_out, I0 =>  inp_feat(62), I1 =>  inp_feat(120), I2 =>  inp_feat(476), I3 =>  inp_feat(277), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_3_L_3_inst : LUT6 generic map(INIT => "1000001100010011000010010010001101001010011111110001011101111111") port map( O =>C_25_S_3_L_3_out, I0 =>  inp_feat(127), I1 =>  inp_feat(67), I2 =>  inp_feat(94), I3 =>  inp_feat(140), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_3_L_4_inst : LUT6 generic map(INIT => "0011011111010000101100011100000001011111110000000111111100000000") port map( O =>C_25_S_3_L_4_out, I0 =>  inp_feat(94), I1 =>  inp_feat(187), I2 =>  inp_feat(389), I3 =>  inp_feat(392), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_3_L_5_inst : LUT6 generic map(INIT => "1111000110001100001001011010000001111100111000001110000010111000") port map( O =>C_25_S_3_L_5_out, I0 =>  inp_feat(472), I1 =>  inp_feat(421), I2 =>  inp_feat(319), I3 =>  inp_feat(503), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_25_S_4_L_0_inst : LUT6 generic map(INIT => "0010101100001101000001010000010100010011111101110011111101111111") port map( O =>C_25_S_4_L_0_out, I0 =>  inp_feat(94), I1 =>  inp_feat(140), I2 =>  inp_feat(67), I3 =>  inp_feat(183), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_4_L_1_inst : LUT6 generic map(INIT => "1111011110001000000000111000100000111111010010000111111100000011") port map( O =>C_25_S_4_L_1_out, I0 =>  inp_feat(389), I1 =>  inp_feat(18), I2 =>  inp_feat(94), I3 =>  inp_feat(279), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_4_L_2_inst : LUT6 generic map(INIT => "0001110110000100001110010000101011110111000000000111111100000000") port map( O =>C_25_S_4_L_2_out, I0 =>  inp_feat(18), I1 =>  inp_feat(94), I2 =>  inp_feat(415), I3 =>  inp_feat(392), I4 =>  inp_feat(275), I5 =>  inp_feat(287)); 
C_25_S_4_L_3_inst : LUT6 generic map(INIT => "0011000110011010011010100010101010000111000110110000111110111011") port map( O =>C_25_S_4_L_3_out, I0 =>  inp_feat(160), I1 =>  inp_feat(354), I2 =>  inp_feat(421), I3 =>  inp_feat(287), I4 =>  inp_feat(169), I5 =>  inp_feat(107)); 
C_25_S_4_L_4_inst : LUT6 generic map(INIT => "1001100011011000110011000101010000000000000010000000000000000000") port map( O =>C_25_S_4_L_4_out, I0 =>  inp_feat(106), I1 =>  inp_feat(292), I2 =>  inp_feat(326), I3 =>  inp_feat(386), I4 =>  inp_feat(363), I5 =>  inp_feat(405)); 
C_25_S_4_L_5_inst : LUT6 generic map(INIT => "0111111111011111100100110000100010011001001110100101001100000000") port map( O =>C_25_S_4_L_5_out, I0 =>  inp_feat(49), I1 =>  inp_feat(421), I2 =>  inp_feat(74), I3 =>  inp_feat(226), I4 =>  inp_feat(307), I5 =>  inp_feat(510)); 
C_25_S_5_L_0_inst : LUT6 generic map(INIT => "0010111001010110110010100000000011110011000101001010101100001010") port map( O =>C_25_S_5_L_0_out, I0 =>  inp_feat(316), I1 =>  inp_feat(167), I2 =>  inp_feat(304), I3 =>  inp_feat(392), I4 =>  inp_feat(473), I5 =>  inp_feat(503)); 
C_25_S_5_L_1_inst : LUT6 generic map(INIT => "0100100110110001000101111111011111011110101010001001000000001001") port map( O =>C_25_S_5_L_1_out, I0 =>  inp_feat(374), I1 =>  inp_feat(354), I2 =>  inp_feat(180), I3 =>  inp_feat(94), I4 =>  inp_feat(20), I5 =>  inp_feat(480)); 
C_25_S_5_L_2_inst : LUT6 generic map(INIT => "1000100100001101000001001111000111101110011011110000001000011111") port map( O =>C_25_S_5_L_2_out, I0 =>  inp_feat(126), I1 =>  inp_feat(507), I2 =>  inp_feat(35), I3 =>  inp_feat(269), I4 =>  inp_feat(299), I5 =>  inp_feat(303)); 
C_25_S_5_L_3_inst : LUT6 generic map(INIT => "0101010101110010000001010001001011101010001010000000000000001000") port map( O =>C_25_S_5_L_3_out, I0 =>  inp_feat(475), I1 =>  inp_feat(163), I2 =>  inp_feat(437), I3 =>  inp_feat(310), I4 =>  inp_feat(145), I5 =>  inp_feat(399)); 
C_25_S_5_L_4_inst : LUT6 generic map(INIT => "1101011001100110000111100010101111011111000001100000001010111111") port map( O =>C_25_S_5_L_4_out, I0 =>  inp_feat(81), I1 =>  inp_feat(421), I2 =>  inp_feat(374), I3 =>  inp_feat(287), I4 =>  inp_feat(127), I5 =>  inp_feat(202)); 
C_25_S_5_L_5_inst : LUT6 generic map(INIT => "0001101100100000100110010000000011111011111110100100000000010011") port map( O =>C_25_S_5_L_5_out, I0 =>  inp_feat(84), I1 =>  inp_feat(441), I2 =>  inp_feat(151), I3 =>  inp_feat(226), I4 =>  inp_feat(307), I5 =>  inp_feat(111)); 
C_26_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111111010000011111111111010001110110010000000") port map( O =>C_26_S_0_L_0_out, I0 =>  inp_feat(167), I1 =>  inp_feat(67), I2 =>  inp_feat(389), I3 =>  inp_feat(421), I4 =>  inp_feat(354), I5 =>  inp_feat(287)); 
C_26_S_0_L_1_inst : LUT6 generic map(INIT => "1110010001111100001111000000000100000001000000010000101100010001") port map( O =>C_26_S_0_L_1_out, I0 =>  inp_feat(399), I1 =>  inp_feat(318), I2 =>  inp_feat(35), I3 =>  inp_feat(127), I4 =>  inp_feat(45), I5 =>  inp_feat(121)); 
C_26_S_0_L_2_inst : LUT6 generic map(INIT => "0010001100001110011000011100100000100001001011110001000011000000") port map( O =>C_26_S_0_L_2_out, I0 =>  inp_feat(335), I1 =>  inp_feat(74), I2 =>  inp_feat(46), I3 =>  inp_feat(279), I4 =>  inp_feat(354), I5 =>  inp_feat(261)); 
C_26_S_0_L_3_inst : LUT6 generic map(INIT => "1011010011101110100010100000100000011000001011001010101000000000") port map( O =>C_26_S_0_L_3_out, I0 =>  inp_feat(354), I1 =>  inp_feat(51), I2 =>  inp_feat(194), I3 =>  inp_feat(127), I4 =>  inp_feat(46), I5 =>  inp_feat(14)); 
C_26_S_0_L_4_inst : LUT6 generic map(INIT => "1100011111110110100110010000011100000001001111110010001000000000") port map( O =>C_26_S_0_L_4_out, I0 =>  inp_feat(386), I1 =>  inp_feat(104), I2 =>  inp_feat(368), I3 =>  inp_feat(45), I4 =>  inp_feat(94), I5 =>  inp_feat(195)); 
C_26_S_0_L_5_inst : LUT6 generic map(INIT => "0011001100100010001101111110111000100001111110111111011101100100") port map( O =>C_26_S_0_L_5_out, I0 =>  inp_feat(403), I1 =>  inp_feat(123), I2 =>  inp_feat(180), I3 =>  inp_feat(448), I4 =>  inp_feat(344), I5 =>  inp_feat(186)); 
C_26_S_1_L_0_inst : LUT6 generic map(INIT => "1110010001111100001111000000000100000001000000010000101100010001") port map( O =>C_26_S_1_L_0_out, I0 =>  inp_feat(399), I1 =>  inp_feat(318), I2 =>  inp_feat(35), I3 =>  inp_feat(127), I4 =>  inp_feat(45), I5 =>  inp_feat(121)); 
C_26_S_1_L_1_inst : LUT6 generic map(INIT => "0010001100001110011000011100100000100001001011110001000011000000") port map( O =>C_26_S_1_L_1_out, I0 =>  inp_feat(335), I1 =>  inp_feat(74), I2 =>  inp_feat(46), I3 =>  inp_feat(279), I4 =>  inp_feat(354), I5 =>  inp_feat(261)); 
C_26_S_1_L_2_inst : LUT6 generic map(INIT => "1011010011101110100010100000100000011000001011001010101000000000") port map( O =>C_26_S_1_L_2_out, I0 =>  inp_feat(354), I1 =>  inp_feat(51), I2 =>  inp_feat(194), I3 =>  inp_feat(127), I4 =>  inp_feat(46), I5 =>  inp_feat(14)); 
C_26_S_1_L_3_inst : LUT6 generic map(INIT => "1100011111110110100110010000011100000001001111110010001000000000") port map( O =>C_26_S_1_L_3_out, I0 =>  inp_feat(386), I1 =>  inp_feat(104), I2 =>  inp_feat(368), I3 =>  inp_feat(45), I4 =>  inp_feat(94), I5 =>  inp_feat(195)); 
C_26_S_1_L_4_inst : LUT6 generic map(INIT => "0011001100100010001101111110111000100001111110111111011101100100") port map( O =>C_26_S_1_L_4_out, I0 =>  inp_feat(403), I1 =>  inp_feat(123), I2 =>  inp_feat(180), I3 =>  inp_feat(448), I4 =>  inp_feat(344), I5 =>  inp_feat(186)); 
C_26_S_1_L_5_inst : LUT6 generic map(INIT => "1010101011100101110101111111000101100111011011100001010010011000") port map( O =>C_26_S_1_L_5_out, I0 =>  inp_feat(17), I1 =>  inp_feat(91), I2 =>  inp_feat(357), I3 =>  inp_feat(102), I4 =>  inp_feat(46), I5 =>  inp_feat(107)); 
C_26_S_2_L_0_inst : LUT6 generic map(INIT => "0000010111101111100111011110111000111011000111000000010011000100") port map( O =>C_26_S_2_L_0_out, I0 =>  inp_feat(334), I1 =>  inp_feat(87), I2 =>  inp_feat(332), I3 =>  inp_feat(292), I4 =>  inp_feat(45), I5 =>  inp_feat(395)); 
C_26_S_2_L_1_inst : LUT6 generic map(INIT => "1110011000011101101000101100100000011010000111110010000011000000") port map( O =>C_26_S_2_L_1_out, I0 =>  inp_feat(503), I1 =>  inp_feat(74), I2 =>  inp_feat(46), I3 =>  inp_feat(279), I4 =>  inp_feat(354), I5 =>  inp_feat(261)); 
C_26_S_2_L_2_inst : LUT6 generic map(INIT => "0011010110011111110101010011110100001101111110100101000011110000") port map( O =>C_26_S_2_L_2_out, I0 =>  inp_feat(92), I1 =>  inp_feat(67), I2 =>  inp_feat(421), I3 =>  inp_feat(279), I4 =>  inp_feat(261), I5 =>  inp_feat(354)); 
C_26_S_2_L_3_inst : LUT6 generic map(INIT => "1111011011001111000001101100111001111111000010111000111001001100") port map( O =>C_26_S_2_L_3_out, I0 =>  inp_feat(323), I1 =>  inp_feat(287), I2 =>  inp_feat(279), I3 =>  inp_feat(18), I4 =>  inp_feat(261), I5 =>  inp_feat(354)); 
C_26_S_2_L_4_inst : LUT6 generic map(INIT => "1111110000100110001101111000111100111110000011000000110000001000") port map( O =>C_26_S_2_L_4_out, I0 =>  inp_feat(67), I1 =>  inp_feat(417), I2 =>  inp_feat(282), I3 =>  inp_feat(107), I4 =>  inp_feat(127), I5 =>  inp_feat(45)); 
C_26_S_2_L_5_inst : LUT6 generic map(INIT => "0101010001011110010001100101110011101110110000001100111011000100") port map( O =>C_26_S_2_L_5_out, I0 =>  inp_feat(138), I1 =>  inp_feat(127), I2 =>  inp_feat(88), I3 =>  inp_feat(452), I4 =>  inp_feat(398), I5 =>  inp_feat(487)); 
C_26_S_3_L_0_inst : LUT6 generic map(INIT => "1111111111001001001001101000100000101111000011110000110000001100") port map( O =>C_26_S_3_L_0_out, I0 =>  inp_feat(67), I1 =>  inp_feat(421), I2 =>  inp_feat(279), I3 =>  inp_feat(18), I4 =>  inp_feat(261), I5 =>  inp_feat(354)); 
C_26_S_3_L_1_inst : LUT6 generic map(INIT => "0100011100010101101010111011001011110111011101010011001000110000") port map( O =>C_26_S_3_L_1_out, I0 =>  inp_feat(70), I1 =>  inp_feat(15), I2 =>  inp_feat(18), I3 =>  inp_feat(140), I4 =>  inp_feat(261), I5 =>  inp_feat(287)); 
C_26_S_3_L_2_inst : LUT6 generic map(INIT => "1111010111001111011100001111010101010010101110100101000010110010") port map( O =>C_26_S_3_L_2_out, I0 =>  inp_feat(31), I1 =>  inp_feat(166), I2 =>  inp_feat(395), I3 =>  inp_feat(321), I4 =>  inp_feat(169), I5 =>  inp_feat(287)); 
C_26_S_3_L_3_inst : LUT6 generic map(INIT => "1000000001100000010000100110001010101100111011001110000011101100") port map( O =>C_26_S_3_L_3_out, I0 =>  inp_feat(45), I1 =>  inp_feat(419), I2 =>  inp_feat(145), I3 =>  inp_feat(159), I4 =>  inp_feat(398), I5 =>  inp_feat(487)); 
C_26_S_3_L_4_inst : LUT6 generic map(INIT => "0100111111000111111001111101111100000000011001101110011111011111") port map( O =>C_26_S_3_L_4_out, I0 =>  inp_feat(374), I1 =>  inp_feat(18), I2 =>  inp_feat(159), I3 =>  inp_feat(398), I4 =>  inp_feat(487), I5 =>  inp_feat(456)); 
C_26_S_3_L_5_inst : LUT6 generic map(INIT => "0111011000011110001101001011011011111110111011100010111011101110") port map( O =>C_26_S_3_L_5_out, I0 =>  inp_feat(368), I1 =>  inp_feat(242), I2 =>  inp_feat(239), I3 =>  inp_feat(389), I4 =>  inp_feat(1), I5 =>  inp_feat(204)); 
C_26_S_4_L_0_inst : LUT6 generic map(INIT => "1100111011001010101011101110110000101010100011101000100001001000") port map( O =>C_26_S_4_L_0_out, I0 =>  inp_feat(503), I1 =>  inp_feat(18), I2 =>  inp_feat(183), I3 =>  inp_feat(249), I4 =>  inp_feat(395), I5 =>  inp_feat(45)); 
C_26_S_4_L_1_inst : LUT6 generic map(INIT => "1110100000110001010110110011001100010000111100110010001000100010") port map( O =>C_26_S_4_L_1_out, I0 =>  inp_feat(67), I1 =>  inp_feat(480), I2 =>  inp_feat(140), I3 =>  inp_feat(183), I4 =>  inp_feat(127), I5 =>  inp_feat(484)); 
C_26_S_4_L_2_inst : LUT6 generic map(INIT => "0000001010100110000000001110000011101111111111100100000011000000") port map( O =>C_26_S_4_L_2_out, I0 =>  inp_feat(492), I1 =>  inp_feat(127), I2 =>  inp_feat(242), I3 =>  inp_feat(305), I4 =>  inp_feat(169), I5 =>  inp_feat(401)); 
C_26_S_4_L_3_inst : LUT6 generic map(INIT => "0110110011011111110111111101111111111101101111111111111111110110") port map( O =>C_26_S_4_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(361), I2 =>  inp_feat(322), I3 =>  inp_feat(392), I4 =>  inp_feat(482), I5 =>  inp_feat(124)); 
C_26_S_4_L_4_inst : LUT6 generic map(INIT => "0000110010101011001010101011111110110011101101101111101111111111") port map( O =>C_26_S_4_L_4_out, I0 =>  inp_feat(395), I1 =>  inp_feat(336), I2 =>  inp_feat(38), I3 =>  inp_feat(55), I4 =>  inp_feat(40), I5 =>  inp_feat(31)); 
C_26_S_4_L_5_inst : LUT6 generic map(INIT => "1111111111100010111111110000110000100010001001101110011100000100") port map( O =>C_26_S_4_L_5_out, I0 =>  inp_feat(140), I1 =>  inp_feat(287), I2 =>  inp_feat(253), I3 =>  inp_feat(94), I4 =>  inp_feat(45), I5 =>  inp_feat(456)); 
C_26_S_5_L_0_inst : LUT6 generic map(INIT => "0000000010110100011011011111000000011111011100011101111111111100") port map( O =>C_26_S_5_L_0_out, I0 =>  inp_feat(44), I1 =>  inp_feat(71), I2 =>  inp_feat(241), I3 =>  inp_feat(251), I4 =>  inp_feat(476), I5 =>  inp_feat(403)); 
C_26_S_5_L_1_inst : LUT6 generic map(INIT => "1111100010111011111000111100000000000010111110111010000000010000") port map( O =>C_26_S_5_L_1_out, I0 =>  inp_feat(503), I1 =>  inp_feat(211), I2 =>  inp_feat(167), I3 =>  inp_feat(249), I4 =>  inp_feat(46), I5 =>  inp_feat(127)); 
C_26_S_5_L_2_inst : LUT6 generic map(INIT => "0001010111100101110101111000110000010000111101001111011110000011") port map( O =>C_26_S_5_L_2_out, I0 =>  inp_feat(438), I1 =>  inp_feat(216), I2 =>  inp_feat(37), I3 =>  inp_feat(70), I4 =>  inp_feat(458), I5 =>  inp_feat(484)); 
C_26_S_5_L_3_inst : LUT6 generic map(INIT => "1110110011110111011001001011100011111010111100100000000011110000") port map( O =>C_26_S_5_L_3_out, I0 =>  inp_feat(183), I1 =>  inp_feat(127), I2 =>  inp_feat(67), I3 =>  inp_feat(123), I4 =>  inp_feat(144), I5 =>  inp_feat(401)); 
C_26_S_5_L_4_inst : LUT6 generic map(INIT => "0010011001111000001001101110100001001100111010001111110011110000") port map( O =>C_26_S_5_L_4_out, I0 =>  inp_feat(94), I1 =>  inp_feat(503), I2 =>  inp_feat(107), I3 =>  inp_feat(304), I4 =>  inp_feat(336), I5 =>  inp_feat(220)); 
C_26_S_5_L_5_inst : LUT6 generic map(INIT => "1010101011101110111111001101111000100000001011110010110011101111") port map( O =>C_26_S_5_L_5_out, I0 =>  inp_feat(503), I1 =>  inp_feat(421), I2 =>  inp_feat(375), I3 =>  inp_feat(93), I4 =>  inp_feat(68), I5 =>  inp_feat(404)); 
C_27_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111111110100011111111111010001110110010000000") port map( O =>C_27_S_0_L_0_out, I0 =>  inp_feat(127), I1 =>  inp_feat(67), I2 =>  inp_feat(389), I3 =>  inp_feat(421), I4 =>  inp_feat(354), I5 =>  inp_feat(287)); 
C_27_S_0_L_1_inst : LUT6 generic map(INIT => "1111111100101011000001101111110000101011100010100000000000110111") port map( O =>C_27_S_0_L_1_out, I0 =>  inp_feat(288), I1 =>  inp_feat(231), I2 =>  inp_feat(320), I3 =>  inp_feat(455), I4 =>  inp_feat(389), I5 =>  inp_feat(169)); 
C_27_S_0_L_2_inst : LUT6 generic map(INIT => "1011000111110111001100111101011100110000001000100010000011000000") port map( O =>C_27_S_0_L_2_out, I0 =>  inp_feat(251), I1 =>  inp_feat(488), I2 =>  inp_feat(220), I3 =>  inp_feat(480), I4 =>  inp_feat(127), I5 =>  inp_feat(46)); 
C_27_S_0_L_3_inst : LUT6 generic map(INIT => "0110000000101011111111011110111011111111110110001111110011110000") port map( O =>C_27_S_0_L_3_out, I0 =>  inp_feat(464), I1 =>  inp_feat(40), I2 =>  inp_feat(148), I3 =>  inp_feat(379), I4 =>  inp_feat(316), I5 =>  inp_feat(123)); 
C_27_S_0_L_4_inst : LUT6 generic map(INIT => "1111111110011011000011111011100001000011000111110000100011111000") port map( O =>C_27_S_0_L_4_out, I0 =>  inp_feat(87), I1 =>  inp_feat(287), I2 =>  inp_feat(245), I3 =>  inp_feat(226), I4 =>  inp_feat(503), I5 =>  inp_feat(18)); 
C_27_S_0_L_5_inst : LUT6 generic map(INIT => "1010010000100011001001101110010011101110111010001110010011101100") port map( O =>C_27_S_0_L_5_out, I0 =>  inp_feat(287), I1 =>  inp_feat(94), I2 =>  inp_feat(67), I3 =>  inp_feat(485), I4 =>  inp_feat(115), I5 =>  inp_feat(155)); 
C_27_S_1_L_0_inst : LUT6 generic map(INIT => "1111111100101011000001101111110000101011100010100000000000110111") port map( O =>C_27_S_1_L_0_out, I0 =>  inp_feat(288), I1 =>  inp_feat(231), I2 =>  inp_feat(320), I3 =>  inp_feat(455), I4 =>  inp_feat(389), I5 =>  inp_feat(169)); 
C_27_S_1_L_1_inst : LUT6 generic map(INIT => "1011000111110111001100111101011100110000001000100010000011000000") port map( O =>C_27_S_1_L_1_out, I0 =>  inp_feat(251), I1 =>  inp_feat(488), I2 =>  inp_feat(220), I3 =>  inp_feat(480), I4 =>  inp_feat(127), I5 =>  inp_feat(46)); 
C_27_S_1_L_2_inst : LUT6 generic map(INIT => "0110000000101011111111011110111011111111110110001111110011110000") port map( O =>C_27_S_1_L_2_out, I0 =>  inp_feat(464), I1 =>  inp_feat(40), I2 =>  inp_feat(148), I3 =>  inp_feat(379), I4 =>  inp_feat(316), I5 =>  inp_feat(123)); 
C_27_S_1_L_3_inst : LUT6 generic map(INIT => "1111111110011011000011111011100001000011000111110000100011111000") port map( O =>C_27_S_1_L_3_out, I0 =>  inp_feat(87), I1 =>  inp_feat(287), I2 =>  inp_feat(245), I3 =>  inp_feat(226), I4 =>  inp_feat(503), I5 =>  inp_feat(18)); 
C_27_S_1_L_4_inst : LUT6 generic map(INIT => "1010010000100011001001101110010011101110111010001110010011101100") port map( O =>C_27_S_1_L_4_out, I0 =>  inp_feat(287), I1 =>  inp_feat(94), I2 =>  inp_feat(67), I3 =>  inp_feat(485), I4 =>  inp_feat(115), I5 =>  inp_feat(155)); 
C_27_S_1_L_5_inst : LUT6 generic map(INIT => "0010001000011111010111100011100011111101011110000011100000101010") port map( O =>C_27_S_1_L_5_out, I0 =>  inp_feat(440), I1 =>  inp_feat(504), I2 =>  inp_feat(488), I3 =>  inp_feat(311), I4 =>  inp_feat(493), I5 =>  inp_feat(445)); 
C_27_S_2_L_0_inst : LUT6 generic map(INIT => "1111000010101100000100101101111110000010111101100100010100001100") port map( O =>C_27_S_2_L_0_out, I0 =>  inp_feat(242), I1 =>  inp_feat(311), I2 =>  inp_feat(194), I3 =>  inp_feat(489), I4 =>  inp_feat(354), I5 =>  inp_feat(261)); 
C_27_S_2_L_1_inst : LUT6 generic map(INIT => "1101100000111010100111000000000001011100001000000010000010000000") port map( O =>C_27_S_2_L_1_out, I0 =>  inp_feat(195), I1 =>  inp_feat(287), I2 =>  inp_feat(94), I3 =>  inp_feat(67), I4 =>  inp_feat(261), I5 =>  inp_feat(374)); 
C_27_S_2_L_2_inst : LUT6 generic map(INIT => "0111001100100010011000111110000011111110110010000111101011100000") port map( O =>C_27_S_2_L_2_out, I0 =>  inp_feat(208), I1 =>  inp_feat(170), I2 =>  inp_feat(130), I3 =>  inp_feat(118), I4 =>  inp_feat(78), I5 =>  inp_feat(284)); 
C_27_S_2_L_3_inst : LUT6 generic map(INIT => "1011110111110111010011001100011111111111011111111111111111110010") port map( O =>C_27_S_2_L_3_out, I0 =>  inp_feat(453), I1 =>  inp_feat(280), I2 =>  inp_feat(207), I3 =>  inp_feat(143), I4 =>  inp_feat(73), I5 =>  inp_feat(155)); 
C_27_S_2_L_4_inst : LUT6 generic map(INIT => "1011010110101111111011110001101000001000001111010000100011001100") port map( O =>C_27_S_2_L_4_out, I0 =>  inp_feat(389), I1 =>  inp_feat(249), I2 =>  inp_feat(92), I3 =>  inp_feat(226), I4 =>  inp_feat(503), I5 =>  inp_feat(18)); 
C_27_S_2_L_5_inst : LUT6 generic map(INIT => "1001100100010111011101001111010000011101000101010000000011110000") port map( O =>C_27_S_2_L_5_out, I0 =>  inp_feat(489), I1 =>  inp_feat(94), I2 =>  inp_feat(287), I3 =>  inp_feat(250), I4 =>  inp_feat(140), I5 =>  inp_feat(167)); 
C_27_S_3_L_0_inst : LUT6 generic map(INIT => "1001111111011100001000010010111011011110111111000010111111111100") port map( O =>C_27_S_3_L_0_out, I0 =>  inp_feat(160), I1 =>  inp_feat(421), I2 =>  inp_feat(212), I3 =>  inp_feat(91), I4 =>  inp_feat(73), I5 =>  inp_feat(155)); 
C_27_S_3_L_1_inst : LUT6 generic map(INIT => "1010100010111000111110101110100000101010001000100001101011111000") port map( O =>C_27_S_3_L_1_out, I0 =>  inp_feat(417), I1 =>  inp_feat(139), I2 =>  inp_feat(347), I3 =>  inp_feat(169), I4 =>  inp_feat(194), I5 =>  inp_feat(121)); 
C_27_S_3_L_2_inst : LUT6 generic map(INIT => "0001101011010100010001000001000001011100111100010001000011000101") port map( O =>C_27_S_3_L_2_out, I0 =>  inp_feat(445), I1 =>  inp_feat(167), I2 =>  inp_feat(311), I3 =>  inp_feat(194), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_27_S_3_L_3_inst : LUT6 generic map(INIT => "0010101100000011011101101101110111111111111011011111111111111110") port map( O =>C_27_S_3_L_3_out, I0 =>  inp_feat(374), I1 =>  inp_feat(404), I2 =>  inp_feat(504), I3 =>  inp_feat(421), I4 =>  inp_feat(73), I5 =>  inp_feat(155)); 
C_27_S_3_L_4_inst : LUT6 generic map(INIT => "1011101111110010111110101110001000101111111100100001000001110000") port map( O =>C_27_S_3_L_4_out, I0 =>  inp_feat(287), I1 =>  inp_feat(418), I2 =>  inp_feat(94), I3 =>  inp_feat(45), I4 =>  inp_feat(65), I5 =>  inp_feat(29)); 
C_27_S_3_L_5_inst : LUT6 generic map(INIT => "0011101111110010111100100010001100011000101100001111101000100000") port map( O =>C_27_S_3_L_5_out, I0 =>  inp_feat(503), I1 =>  inp_feat(289), I2 =>  inp_feat(18), I3 =>  inp_feat(395), I4 =>  inp_feat(45), I5 =>  inp_feat(448)); 
C_27_S_4_L_0_inst : LUT6 generic map(INIT => "1000101100000111000000111011111101010010100111010000001110011011") port map( O =>C_27_S_4_L_0_out, I0 =>  inp_feat(354), I1 =>  inp_feat(215), I2 =>  inp_feat(456), I3 =>  inp_feat(489), I4 =>  inp_feat(503), I5 =>  inp_feat(18)); 
C_27_S_4_L_1_inst : LUT6 generic map(INIT => "1010101000111111011111111010000011111011000010110001100000100000") port map( O =>C_27_S_4_L_1_out, I0 =>  inp_feat(395), I1 =>  inp_feat(282), I2 =>  inp_feat(250), I3 =>  inp_feat(127), I4 =>  inp_feat(31), I5 =>  inp_feat(220)); 
C_27_S_4_L_2_inst : LUT6 generic map(INIT => "0001010000011101111110100011100011111101111110111100000000000000") port map( O =>C_27_S_4_L_2_out, I0 =>  inp_feat(446), I1 =>  inp_feat(450), I2 =>  inp_feat(405), I3 =>  inp_feat(493), I4 =>  inp_feat(390), I5 =>  inp_feat(358)); 
C_27_S_4_L_3_inst : LUT6 generic map(INIT => "1011110001101111110011001111101110010100010111110100110011011000") port map( O =>C_27_S_4_L_3_out, I0 =>  inp_feat(244), I1 =>  inp_feat(420), I2 =>  inp_feat(48), I3 =>  inp_feat(389), I4 =>  inp_feat(114), I5 =>  inp_feat(448)); 
C_27_S_4_L_4_inst : LUT6 generic map(INIT => "1101110110111100101000101101000000010111101111000000000001100010") port map( O =>C_27_S_4_L_4_out, I0 =>  inp_feat(427), I1 =>  inp_feat(186), I2 =>  inp_feat(311), I3 =>  inp_feat(194), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_27_S_4_L_5_inst : LUT6 generic map(INIT => "1110011001111010111001111111001001111010000010000111001011101111") port map( O =>C_27_S_4_L_5_out, I0 =>  inp_feat(153), I1 =>  inp_feat(212), I2 =>  inp_feat(490), I3 =>  inp_feat(385), I4 =>  inp_feat(261), I5 =>  inp_feat(374)); 
C_27_S_5_L_0_inst : LUT6 generic map(INIT => "0001100110100010000001111111101111111111111111001010111111111110") port map( O =>C_27_S_5_L_0_out, I0 =>  inp_feat(208), I1 =>  inp_feat(45), I2 =>  inp_feat(6), I3 =>  inp_feat(212), I4 =>  inp_feat(73), I5 =>  inp_feat(155)); 
C_27_S_5_L_1_inst : LUT6 generic map(INIT => "1100001011001111110111111000011100000111101111111111111100111111") port map( O =>C_27_S_5_L_1_out, I0 =>  inp_feat(250), I1 =>  inp_feat(101), I2 =>  inp_feat(480), I3 =>  inp_feat(118), I4 =>  inp_feat(263), I5 =>  inp_feat(37)); 
C_27_S_5_L_2_inst : LUT6 generic map(INIT => "0111111100011101101011011111110111011100010010000100010001000000") port map( O =>C_27_S_5_L_2_out, I0 =>  inp_feat(257), I1 =>  inp_feat(45), I2 =>  inp_feat(172), I3 =>  inp_feat(127), I4 =>  inp_feat(288), I5 =>  inp_feat(220)); 
C_27_S_5_L_3_inst : LUT6 generic map(INIT => "1011100011111111111100101111111111110010111111110010001011111011") port map( O =>C_27_S_5_L_3_out, I0 =>  inp_feat(171), I1 =>  inp_feat(445), I2 =>  inp_feat(291), I3 =>  inp_feat(308), I4 =>  inp_feat(429), I5 =>  inp_feat(106)); 
C_27_S_5_L_4_inst : LUT6 generic map(INIT => "0111001000000010100010000110001011111111101000101110101101100010") port map( O =>C_27_S_5_L_4_out, I0 =>  inp_feat(169), I1 =>  inp_feat(59), I2 =>  inp_feat(46), I3 =>  inp_feat(354), I4 =>  inp_feat(189), I5 =>  inp_feat(295)); 
C_27_S_5_L_5_inst : LUT6 generic map(INIT => "0000010010000110111011000000000011111110111011001100010010000100") port map( O =>C_27_S_5_L_5_out, I0 =>  inp_feat(287), I1 =>  inp_feat(484), I2 =>  inp_feat(420), I3 =>  inp_feat(265), I4 =>  inp_feat(370), I5 =>  inp_feat(174)); 
C_28_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000010000011100000000000111110000011101111111") port map( O =>C_28_S_0_L_0_out, I0 =>  inp_feat(18), I1 =>  inp_feat(67), I2 =>  inp_feat(389), I3 =>  inp_feat(421), I4 =>  inp_feat(354), I5 =>  inp_feat(287)); 
C_28_S_0_L_1_inst : LUT6 generic map(INIT => "0000000101000100111001100000110011101111100011111110111110001110") port map( O =>C_28_S_0_L_1_out, I0 =>  inp_feat(472), I1 =>  inp_feat(182), I2 =>  inp_feat(493), I3 =>  inp_feat(1), I4 =>  inp_feat(127), I5 =>  inp_feat(497)); 
C_28_S_0_L_2_inst : LUT6 generic map(INIT => "0100100110111101010000100111000100111010111100010111111111110111") port map( O =>C_28_S_0_L_2_out, I0 =>  inp_feat(389), I1 =>  inp_feat(354), I2 =>  inp_feat(455), I3 =>  inp_feat(46), I4 =>  inp_feat(37), I5 =>  inp_feat(374)); 
C_28_S_0_L_3_inst : LUT6 generic map(INIT => "0101100111111000010101011111100011011110111101001001000011101000") port map( O =>C_28_S_0_L_3_out, I0 =>  inp_feat(470), I1 =>  inp_feat(157), I2 =>  inp_feat(101), I3 =>  inp_feat(503), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_28_S_0_L_4_inst : LUT6 generic map(INIT => "0101011101000001111100111001000110110111000000110011111100100111") port map( O =>C_28_S_0_L_4_out, I0 =>  inp_feat(67), I1 =>  inp_feat(140), I2 =>  inp_feat(287), I3 =>  inp_feat(111), I4 =>  inp_feat(354), I5 =>  inp_feat(49)); 
C_28_S_0_L_5_inst : LUT6 generic map(INIT => "1010100000010010111001110000000010110011000010001111111100000010") port map( O =>C_28_S_0_L_5_out, I0 =>  inp_feat(25), I1 =>  inp_feat(67), I2 =>  inp_feat(3), I3 =>  inp_feat(478), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_28_S_1_L_0_inst : LUT6 generic map(INIT => "0000000101000100111001100000110011101111100011111110111110001110") port map( O =>C_28_S_1_L_0_out, I0 =>  inp_feat(472), I1 =>  inp_feat(182), I2 =>  inp_feat(493), I3 =>  inp_feat(1), I4 =>  inp_feat(127), I5 =>  inp_feat(497)); 
C_28_S_1_L_1_inst : LUT6 generic map(INIT => "0100100110111101010000100111000100111010111100010111111111110111") port map( O =>C_28_S_1_L_1_out, I0 =>  inp_feat(389), I1 =>  inp_feat(354), I2 =>  inp_feat(455), I3 =>  inp_feat(46), I4 =>  inp_feat(37), I5 =>  inp_feat(374)); 
C_28_S_1_L_2_inst : LUT6 generic map(INIT => "0101100111111000010101011111100011011110111101001001000011101000") port map( O =>C_28_S_1_L_2_out, I0 =>  inp_feat(470), I1 =>  inp_feat(157), I2 =>  inp_feat(101), I3 =>  inp_feat(503), I4 =>  inp_feat(261), I5 =>  inp_feat(107)); 
C_28_S_1_L_3_inst : LUT6 generic map(INIT => "0101011101000001111100111001000110110111000000110011111100100111") port map( O =>C_28_S_1_L_3_out, I0 =>  inp_feat(67), I1 =>  inp_feat(140), I2 =>  inp_feat(287), I3 =>  inp_feat(111), I4 =>  inp_feat(354), I5 =>  inp_feat(49)); 
C_28_S_1_L_4_inst : LUT6 generic map(INIT => "1010100000010010111001110000000010110011000010001111111100000010") port map( O =>C_28_S_1_L_4_out, I0 =>  inp_feat(25), I1 =>  inp_feat(67), I2 =>  inp_feat(3), I3 =>  inp_feat(478), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_28_S_1_L_5_inst : LUT6 generic map(INIT => "0011101010000010000001011100000011111010000000000000000000000000") port map( O =>C_28_S_1_L_5_out, I0 =>  inp_feat(282), I1 =>  inp_feat(94), I2 =>  inp_feat(473), I3 =>  inp_feat(371), I4 =>  inp_feat(326), I5 =>  inp_feat(109)); 
C_28_S_2_L_0_inst : LUT6 generic map(INIT => "0100011110101111000000110101111111000001000001011111111111111111") port map( O =>C_28_S_2_L_0_out, I0 =>  inp_feat(94), I1 =>  inp_feat(20), I2 =>  inp_feat(37), I3 =>  inp_feat(374), I4 =>  inp_feat(287), I5 =>  inp_feat(275)); 
C_28_S_2_L_1_inst : LUT6 generic map(INIT => "1100101100101111101010111111101100100010000110010000000000000000") port map( O =>C_28_S_2_L_1_out, I0 =>  inp_feat(48), I1 =>  inp_feat(158), I2 =>  inp_feat(110), I3 =>  inp_feat(258), I4 =>  inp_feat(443), I5 =>  inp_feat(478)); 
C_28_S_2_L_2_inst : LUT6 generic map(INIT => "0110001001010111000000001101111110001111000001010001011110111111") port map( O =>C_28_S_2_L_2_out, I0 =>  inp_feat(127), I1 =>  inp_feat(67), I2 =>  inp_feat(94), I3 =>  inp_feat(374), I4 =>  inp_feat(287), I5 =>  inp_feat(49)); 
C_28_S_2_L_3_inst : LUT6 generic map(INIT => "0000001000011111000000100000110011100001000111111111110100000000") port map( O =>C_28_S_2_L_3_out, I0 =>  inp_feat(395), I1 =>  inp_feat(231), I2 =>  inp_feat(189), I3 =>  inp_feat(55), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_28_S_2_L_4_inst : LUT6 generic map(INIT => "0101010111011101101111011100110111111011000000001010001000000010") port map( O =>C_28_S_2_L_4_out, I0 =>  inp_feat(127), I1 =>  inp_feat(318), I2 =>  inp_feat(107), I3 =>  inp_feat(183), I4 =>  inp_feat(114), I5 =>  inp_feat(388)); 
C_28_S_2_L_5_inst : LUT6 generic map(INIT => "1111110110101100101001000010010000000000100100001001100000000100") port map( O =>C_28_S_2_L_5_out, I0 =>  inp_feat(215), I1 =>  inp_feat(51), I2 =>  inp_feat(263), I3 =>  inp_feat(109), I4 =>  inp_feat(108), I5 =>  inp_feat(391)); 
C_28_S_3_L_0_inst : LUT6 generic map(INIT => "0111010001010010110100110000000011110111000100111111110100001000") port map( O =>C_28_S_3_L_0_out, I0 =>  inp_feat(18), I1 =>  inp_feat(189), I2 =>  inp_feat(219), I3 =>  inp_feat(1), I4 =>  inp_feat(121), I5 =>  inp_feat(110)); 
C_28_S_3_L_1_inst : LUT6 generic map(INIT => "0000000100110000110100100000010010111000001001001000111000001000") port map( O =>C_28_S_3_L_1_out, I0 =>  inp_feat(22), I1 =>  inp_feat(48), I2 =>  inp_feat(287), I3 =>  inp_feat(232), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_28_S_3_L_2_inst : LUT6 generic map(INIT => "0101001001011111010100101110011111111010000010110000001000000010") port map( O =>C_28_S_3_L_2_out, I0 =>  inp_feat(283), I1 =>  inp_feat(94), I2 =>  inp_feat(287), I3 =>  inp_feat(275), I4 =>  inp_feat(379), I5 =>  inp_feat(401)); 
C_28_S_3_L_3_inst : LUT6 generic map(INIT => "1011100100010011000101010001111111010010110100100000101011001010") port map( O =>C_28_S_3_L_3_out, I0 =>  inp_feat(503), I1 =>  inp_feat(183), I2 =>  inp_feat(203), I3 =>  inp_feat(114), I4 =>  inp_feat(164), I5 =>  inp_feat(273)); 
C_28_S_3_L_4_inst : LUT6 generic map(INIT => "0010001101111001000010101101100001010010110100101100001011110000") port map( O =>C_28_S_3_L_4_out, I0 =>  inp_feat(18), I1 =>  inp_feat(318), I2 =>  inp_feat(186), I3 =>  inp_feat(503), I4 =>  inp_feat(323), I5 =>  inp_feat(29)); 
C_28_S_3_L_5_inst : LUT6 generic map(INIT => "1001000110110000000010100000010011111000101001001000111000001000") port map( O =>C_28_S_3_L_5_out, I0 =>  inp_feat(22), I1 =>  inp_feat(48), I2 =>  inp_feat(287), I3 =>  inp_feat(232), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_28_S_4_L_0_inst : LUT6 generic map(INIT => "0000000010110000101000001110000011101010000010001010100010101010") port map( O =>C_28_S_4_L_0_out, I0 =>  inp_feat(445), I1 =>  inp_feat(507), I2 =>  inp_feat(306), I3 =>  inp_feat(503), I4 =>  inp_feat(37), I5 =>  inp_feat(46)); 
C_28_S_4_L_1_inst : LUT6 generic map(INIT => "1010011100111001001000000000000110111111110101001000101100000000") port map( O =>C_28_S_4_L_1_out, I0 =>  inp_feat(101), I1 =>  inp_feat(59), I2 =>  inp_feat(105), I3 =>  inp_feat(251), I4 =>  inp_feat(422), I5 =>  inp_feat(461)); 
C_28_S_4_L_2_inst : LUT6 generic map(INIT => "0000000100111101010101100100001011101000011100000000111011100000") port map( O =>C_28_S_4_L_2_out, I0 =>  inp_feat(108), I1 =>  inp_feat(292), I2 =>  inp_feat(288), I3 =>  inp_feat(277), I4 =>  inp_feat(441), I5 =>  inp_feat(471)); 
C_28_S_4_L_3_inst : LUT6 generic map(INIT => "0100110100101000101011100000001010000111100000001010101000000000") port map( O =>C_28_S_4_L_3_out, I0 =>  inp_feat(392), I1 =>  inp_feat(473), I2 =>  inp_feat(120), I3 =>  inp_feat(289), I4 =>  inp_feat(94), I5 =>  inp_feat(50)); 
C_28_S_4_L_4_inst : LUT6 generic map(INIT => "0101001011010100110001010101111110000100100000000000000000000001") port map( O =>C_28_S_4_L_4_out, I0 =>  inp_feat(374), I1 =>  inp_feat(490), I2 =>  inp_feat(212), I3 =>  inp_feat(114), I4 =>  inp_feat(11), I5 =>  inp_feat(56)); 
C_28_S_4_L_5_inst : LUT6 generic map(INIT => "1011000011001000100100001100100000000010010000001010000011000000") port map( O =>C_28_S_4_L_5_out, I0 =>  inp_feat(422), I1 =>  inp_feat(176), I2 =>  inp_feat(4), I3 =>  inp_feat(225), I4 =>  inp_feat(215), I5 =>  inp_feat(199)); 
C_28_S_5_L_0_inst : LUT6 generic map(INIT => "0110000111011100000000001001000001000001100000001100100010001010") port map( O =>C_28_S_5_L_0_out, I0 =>  inp_feat(403), I1 =>  inp_feat(138), I2 =>  inp_feat(510), I3 =>  inp_feat(313), I4 =>  inp_feat(330), I5 =>  inp_feat(56)); 
C_28_S_5_L_1_inst : LUT6 generic map(INIT => "0001001010100000101100101011101111001100101000101011001011111010") port map( O =>C_28_S_5_L_1_out, I0 =>  inp_feat(13), I1 =>  inp_feat(503), I2 =>  inp_feat(315), I3 =>  inp_feat(94), I4 =>  inp_feat(20), I5 =>  inp_feat(294)); 
C_28_S_5_L_2_inst : LUT6 generic map(INIT => "1101110110100010011011010010001000010010011000101010110110100010") port map( O =>C_28_S_5_L_2_out, I0 =>  inp_feat(199), I1 =>  inp_feat(287), I2 =>  inp_feat(431), I3 =>  inp_feat(275), I4 =>  inp_feat(323), I5 =>  inp_feat(29)); 
C_28_S_5_L_3_inst : LUT6 generic map(INIT => "0000000110000000001010100000011011000000100000000000100000011000") port map( O =>C_28_S_5_L_3_out, I0 =>  inp_feat(454), I1 =>  inp_feat(207), I2 =>  inp_feat(68), I3 =>  inp_feat(57), I4 =>  inp_feat(83), I5 =>  inp_feat(9)); 
C_28_S_5_L_4_inst : LUT6 generic map(INIT => "1110010001001000110011011000000011101100000010001101110100000100") port map( O =>C_28_S_5_L_4_out, I0 =>  inp_feat(287), I1 =>  inp_feat(123), I2 =>  inp_feat(473), I3 =>  inp_feat(257), I4 =>  inp_feat(195), I5 =>  inp_feat(461)); 
C_28_S_5_L_5_inst : LUT6 generic map(INIT => "0001000011010010000001010000001010100101000001001101111100000101") port map( O =>C_28_S_5_L_5_out, I0 =>  inp_feat(389), I1 =>  inp_feat(84), I2 =>  inp_feat(20), I3 =>  inp_feat(151), I4 =>  inp_feat(419), I5 =>  inp_feat(45)); 
C_29_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000000001011100000000000101110001011101111111") port map( O =>C_29_S_0_L_0_out, I0 =>  inp_feat(18), I1 =>  inp_feat(127), I2 =>  inp_feat(389), I3 =>  inp_feat(421), I4 =>  inp_feat(354), I5 =>  inp_feat(287)); 
C_29_S_0_L_1_inst : LUT6 generic map(INIT => "0000000011011000000000001000000010100000111100010000000000000000") port map( O =>C_29_S_0_L_1_out, I0 =>  inp_feat(80), I1 =>  inp_feat(162), I2 =>  inp_feat(449), I3 =>  inp_feat(497), I4 =>  inp_feat(15), I5 =>  inp_feat(121)); 
C_29_S_0_L_2_inst : LUT6 generic map(INIT => "0001000100111101111100000101111110011101101111110011111101111111") port map( O =>C_29_S_0_L_2_out, I0 =>  inp_feat(503), I1 =>  inp_feat(18), I2 =>  inp_feat(287), I3 =>  inp_feat(46), I4 =>  inp_feat(417), I5 =>  inp_feat(356)); 
C_29_S_0_L_3_inst : LUT6 generic map(INIT => "0000011010100010110001000100000000000010000000100001010000000000") port map( O =>C_29_S_0_L_3_out, I0 =>  inp_feat(186), I1 =>  inp_feat(37), I2 =>  inp_feat(287), I3 =>  inp_feat(354), I4 =>  inp_feat(199), I5 =>  inp_feat(282)); 
C_29_S_0_L_4_inst : LUT6 generic map(INIT => "1000101110110100000010011101110000000000001000000000000000000100") port map( O =>C_29_S_0_L_4_out, I0 =>  inp_feat(480), I1 =>  inp_feat(339), I2 =>  inp_feat(168), I3 =>  inp_feat(325), I4 =>  inp_feat(136), I5 =>  inp_feat(15)); 
C_29_S_0_L_5_inst : LUT6 generic map(INIT => "1101100101111000110000000000100001010100000000000000000000000000") port map( O =>C_29_S_0_L_5_out, I0 =>  inp_feat(261), I1 =>  inp_feat(117), I2 =>  inp_feat(40), I3 =>  inp_feat(448), I4 =>  inp_feat(81), I5 =>  inp_feat(246)); 
C_29_S_1_L_0_inst : LUT6 generic map(INIT => "0000000011011000000000001000000010100000111100010000000000000000") port map( O =>C_29_S_1_L_0_out, I0 =>  inp_feat(80), I1 =>  inp_feat(162), I2 =>  inp_feat(449), I3 =>  inp_feat(497), I4 =>  inp_feat(15), I5 =>  inp_feat(121)); 
C_29_S_1_L_1_inst : LUT6 generic map(INIT => "0001000100111101111100000101111110011101101111110011111101111111") port map( O =>C_29_S_1_L_1_out, I0 =>  inp_feat(503), I1 =>  inp_feat(18), I2 =>  inp_feat(287), I3 =>  inp_feat(46), I4 =>  inp_feat(417), I5 =>  inp_feat(356)); 
C_29_S_1_L_2_inst : LUT6 generic map(INIT => "0000011010100010110001000100000000000010000000100001010000000000") port map( O =>C_29_S_1_L_2_out, I0 =>  inp_feat(186), I1 =>  inp_feat(37), I2 =>  inp_feat(287), I3 =>  inp_feat(354), I4 =>  inp_feat(199), I5 =>  inp_feat(282)); 
C_29_S_1_L_3_inst : LUT6 generic map(INIT => "1000101110110100000010011101110000000000001000000000000000000100") port map( O =>C_29_S_1_L_3_out, I0 =>  inp_feat(480), I1 =>  inp_feat(339), I2 =>  inp_feat(168), I3 =>  inp_feat(325), I4 =>  inp_feat(136), I5 =>  inp_feat(15)); 
C_29_S_1_L_4_inst : LUT6 generic map(INIT => "1101100101111000110000000000100001010100000000000000000000000000") port map( O =>C_29_S_1_L_4_out, I0 =>  inp_feat(261), I1 =>  inp_feat(117), I2 =>  inp_feat(40), I3 =>  inp_feat(448), I4 =>  inp_feat(81), I5 =>  inp_feat(246)); 
C_29_S_1_L_5_inst : LUT6 generic map(INIT => "0000001001100001110011011101100000000000000000000000000000001000") port map( O =>C_29_S_1_L_5_out, I0 =>  inp_feat(160), I1 =>  inp_feat(453), I2 =>  inp_feat(168), I3 =>  inp_feat(325), I4 =>  inp_feat(136), I5 =>  inp_feat(15)); 
C_29_S_2_L_0_inst : LUT6 generic map(INIT => "0011001000010010000001010100011000000000000000000000000100100000") port map( O =>C_29_S_2_L_0_out, I0 =>  inp_feat(7), I1 =>  inp_feat(325), I2 =>  inp_feat(445), I3 =>  inp_feat(168), I4 =>  inp_feat(199), I5 =>  inp_feat(15)); 
C_29_S_2_L_1_inst : LUT6 generic map(INIT => "1111011110000010101010001111001000000000000000000001000000000010") port map( O =>C_29_S_2_L_1_out, I0 =>  inp_feat(389), I1 =>  inp_feat(72), I2 =>  inp_feat(228), I3 =>  inp_feat(168), I4 =>  inp_feat(199), I5 =>  inp_feat(15)); 
C_29_S_2_L_2_inst : LUT6 generic map(INIT => "0000010100010111000101110111111100000001000101110000000110001111") port map( O =>C_29_S_2_L_2_out, I0 =>  inp_feat(67), I1 =>  inp_feat(46), I2 =>  inp_feat(261), I3 =>  inp_feat(167), I4 =>  inp_feat(107), I5 =>  inp_feat(98)); 
C_29_S_2_L_3_inst : LUT6 generic map(INIT => "1011000110010011000101010111111100000000010101110000000110010111") port map( O =>C_29_S_2_L_3_out, I0 =>  inp_feat(503), I1 =>  inp_feat(46), I2 =>  inp_feat(261), I3 =>  inp_feat(167), I4 =>  inp_feat(107), I5 =>  inp_feat(98)); 
C_29_S_2_L_4_inst : LUT6 generic map(INIT => "0000100011001101110011001100110100000000000001000000110001001101") port map( O =>C_29_S_2_L_4_out, I0 =>  inp_feat(287), I1 =>  inp_feat(257), I2 =>  inp_feat(167), I3 =>  inp_feat(503), I4 =>  inp_feat(107), I5 =>  inp_feat(312)); 
C_29_S_2_L_5_inst : LUT6 generic map(INIT => "1010010010001100110011000100110100000100000011000100010011001101") port map( O =>C_29_S_2_L_5_out, I0 =>  inp_feat(374), I1 =>  inp_feat(480), I2 =>  inp_feat(37), I3 =>  inp_feat(503), I4 =>  inp_feat(107), I5 =>  inp_feat(312)); 
C_29_S_3_L_0_inst : LUT6 generic map(INIT => "0001001101000011001101110000000100000001000000000000111110000001") port map( O =>C_29_S_3_L_0_out, I0 =>  inp_feat(37), I1 =>  inp_feat(67), I2 =>  inp_feat(261), I3 =>  inp_feat(208), I4 =>  inp_feat(107), I5 =>  inp_feat(98)); 
C_29_S_3_L_1_inst : LUT6 generic map(INIT => "1110111000011100101011000010000000100000000000000010000000100100") port map( O =>C_29_S_3_L_1_out, I0 =>  inp_feat(480), I1 =>  inp_feat(503), I2 =>  inp_feat(168), I3 =>  inp_feat(208), I4 =>  inp_feat(107), I5 =>  inp_feat(98)); 
C_29_S_3_L_2_inst : LUT6 generic map(INIT => "1000101100001000000111110000111100000000000001000000000001000010") port map( O =>C_29_S_3_L_2_out, I0 =>  inp_feat(410), I1 =>  inp_feat(31), I2 =>  inp_feat(281), I3 =>  inp_feat(408), I4 =>  inp_feat(0), I5 =>  inp_feat(387)); 
C_29_S_3_L_3_inst : LUT6 generic map(INIT => "0011000001100000001010001101010100000000010000001111000001000000") port map( O =>C_29_S_3_L_3_out, I0 =>  inp_feat(389), I1 =>  inp_feat(458), I2 =>  inp_feat(448), I3 =>  inp_feat(45), I4 =>  inp_feat(261), I5 =>  inp_feat(246)); 
C_29_S_3_L_4_inst : LUT6 generic map(INIT => "1100011000011000111011000000000000000000000000000100000000100000") port map( O =>C_29_S_3_L_4_out, I0 =>  inp_feat(45), I1 =>  inp_feat(458), I2 =>  inp_feat(448), I3 =>  inp_feat(332), I4 =>  inp_feat(261), I5 =>  inp_feat(246)); 
C_29_S_3_L_5_inst : LUT6 generic map(INIT => "0000000010000000011111110100010000000000000000001000010100001100") port map( O =>C_29_S_3_L_5_out, I0 =>  inp_feat(226), I1 =>  inp_feat(233), I2 =>  inp_feat(418), I3 =>  inp_feat(493), I4 =>  inp_feat(199), I5 =>  inp_feat(471)); 
C_29_S_4_L_0_inst : LUT6 generic map(INIT => "0010100110110000000100000001010000111000011101110000100000100001") port map( O =>C_29_S_4_L_0_out, I0 =>  inp_feat(464), I1 =>  inp_feat(86), I2 =>  inp_feat(275), I3 =>  inp_feat(336), I4 =>  inp_feat(217), I5 =>  inp_feat(281)); 
C_29_S_4_L_1_inst : LUT6 generic map(INIT => "1110100011001111010101011100000101001000001010000000000001000000") port map( O =>C_29_S_4_L_1_out, I0 =>  inp_feat(421), I1 =>  inp_feat(448), I2 =>  inp_feat(335), I3 =>  inp_feat(78), I4 =>  inp_feat(451), I5 =>  inp_feat(84)); 
C_29_S_4_L_2_inst : LUT6 generic map(INIT => "0001011101000111001000110000011100100000001001000000000000000000") port map( O =>C_29_S_4_L_2_out, I0 =>  inp_feat(140), I1 =>  inp_feat(261), I2 =>  inp_feat(287), I3 =>  inp_feat(506), I4 =>  inp_feat(234), I5 =>  inp_feat(209)); 
C_29_S_4_L_3_inst : LUT6 generic map(INIT => "1010010000110010101000000000000000000010000010000000000000000000") port map( O =>C_29_S_4_L_3_out, I0 =>  inp_feat(454), I1 =>  inp_feat(479), I2 =>  inp_feat(79), I3 =>  inp_feat(506), I4 =>  inp_feat(234), I5 =>  inp_feat(209)); 
C_29_S_4_L_4_inst : LUT6 generic map(INIT => "0010000000000000001000100000111000101001000011010001110010001100") port map( O =>C_29_S_4_L_4_out, I0 =>  inp_feat(359), I1 =>  inp_feat(185), I2 =>  inp_feat(319), I3 =>  inp_feat(384), I4 =>  inp_feat(117), I5 =>  inp_feat(474)); 
C_29_S_4_L_5_inst : LUT6 generic map(INIT => "1001110100001000000000000000100010011000100010001000000010001000") port map( O =>C_29_S_4_L_5_out, I0 =>  inp_feat(381), I1 =>  inp_feat(448), I2 =>  inp_feat(344), I3 =>  inp_feat(177), I4 =>  inp_feat(282), I5 =>  inp_feat(403)); 
C_29_S_5_L_0_inst : LUT6 generic map(INIT => "0101110001010011000000110000000011010000000000001000111001011000") port map( O =>C_29_S_5_L_0_out, I0 =>  inp_feat(261), I1 =>  inp_feat(278), I2 =>  inp_feat(143), I3 =>  inp_feat(359), I4 =>  inp_feat(319), I5 =>  inp_feat(281)); 
C_29_S_5_L_1_inst : LUT6 generic map(INIT => "1011111111010101100100110000001100010111000101110000001110000001") port map( O =>C_29_S_5_L_1_out, I0 =>  inp_feat(475), I1 =>  inp_feat(127), I2 =>  inp_feat(389), I3 =>  inp_feat(404), I4 =>  inp_feat(268), I5 =>  inp_feat(246)); 
C_29_S_5_L_2_inst : LUT6 generic map(INIT => "0101000100000000110110110001100111010000100011000001000010001001") port map( O =>C_29_S_5_L_2_out, I0 =>  inp_feat(20), I1 =>  inp_feat(354), I2 =>  inp_feat(135), I3 =>  inp_feat(306), I4 =>  inp_feat(117), I5 =>  inp_feat(489)); 
C_29_S_5_L_3_inst : LUT6 generic map(INIT => "0000000100000111000010100000000011010010100000000000000000000000") port map( O =>C_29_S_5_L_3_out, I0 =>  inp_feat(467), I1 =>  inp_feat(276), I2 =>  inp_feat(4), I3 =>  inp_feat(115), I4 =>  inp_feat(387), I5 =>  inp_feat(43)); 
C_29_S_5_L_4_inst : LUT6 generic map(INIT => "1110100010000001000000010010111100100000000000000000000000000000") port map( O =>C_29_S_5_L_4_out, I0 =>  inp_feat(174), I1 =>  inp_feat(291), I2 =>  inp_feat(96), I3 =>  inp_feat(91), I4 =>  inp_feat(257), I5 =>  inp_feat(387)); 
C_29_S_5_L_5_inst : LUT6 generic map(INIT => "0000000010110100000000000101100011100000101100100000000000000000") port map( O =>C_29_S_5_L_5_out, I0 =>  inp_feat(373), I1 =>  inp_feat(37), I2 =>  inp_feat(41), I3 =>  inp_feat(72), I4 =>  inp_feat(15), I5 =>  inp_feat(374)); 
C_30_S_0_L_0_inst : LUT6 generic map(INIT => "0000000100000001000001010011111100010101000011110001011111111111") port map( O =>C_30_S_0_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(500), I2 =>  inp_feat(307), I3 =>  inp_feat(324), I4 =>  inp_feat(245), I5 =>  inp_feat(424)); 
C_30_S_0_L_1_inst : LUT6 generic map(INIT => "0000011011101101011101111111111110001111111111111111111101111111") port map( O =>C_30_S_0_L_1_out, I0 =>  inp_feat(81), I1 =>  inp_feat(93), I2 =>  inp_feat(210), I3 =>  inp_feat(321), I4 =>  inp_feat(17), I5 =>  inp_feat(489)); 
C_30_S_0_L_2_inst : LUT6 generic map(INIT => "0010100010100000111010101011000111111010101100101011000011111011") port map( O =>C_30_S_0_L_2_out, I0 =>  inp_feat(104), I1 =>  inp_feat(132), I2 =>  inp_feat(292), I3 =>  inp_feat(166), I4 =>  inp_feat(82), I5 =>  inp_feat(255)); 
C_30_S_0_L_3_inst : LUT6 generic map(INIT => "1101110001110101110101000100010001000000000010000000000000000000") port map( O =>C_30_S_0_L_3_out, I0 =>  inp_feat(306), I1 =>  inp_feat(190), I2 =>  inp_feat(94), I3 =>  inp_feat(389), I4 =>  inp_feat(157), I5 =>  inp_feat(221)); 
C_30_S_0_L_4_inst : LUT6 generic map(INIT => "1000010010111100010011001110110000000000000000000000010011111010") port map( O =>C_30_S_0_L_4_out, I0 =>  inp_feat(81), I1 =>  inp_feat(153), I2 =>  inp_feat(65), I3 =>  inp_feat(224), I4 =>  inp_feat(360), I5 =>  inp_feat(84)); 
C_30_S_0_L_5_inst : LUT6 generic map(INIT => "0001000110100010101010011010001000000000001000000110000000100111") port map( O =>C_30_S_0_L_5_out, I0 =>  inp_feat(217), I1 =>  inp_feat(17), I2 =>  inp_feat(292), I3 =>  inp_feat(407), I4 =>  inp_feat(4), I5 =>  inp_feat(75)); 
C_30_S_1_L_0_inst : LUT6 generic map(INIT => "0000011011101101011101111111111110001111111111111111111101111111") port map( O =>C_30_S_1_L_0_out, I0 =>  inp_feat(81), I1 =>  inp_feat(93), I2 =>  inp_feat(210), I3 =>  inp_feat(321), I4 =>  inp_feat(17), I5 =>  inp_feat(489)); 
C_30_S_1_L_1_inst : LUT6 generic map(INIT => "0010100010100000111010101011000111111010101100101011000011111011") port map( O =>C_30_S_1_L_1_out, I0 =>  inp_feat(104), I1 =>  inp_feat(132), I2 =>  inp_feat(292), I3 =>  inp_feat(166), I4 =>  inp_feat(82), I5 =>  inp_feat(255)); 
C_30_S_1_L_2_inst : LUT6 generic map(INIT => "1101110001110101110101000100010001000000000010000000000000000000") port map( O =>C_30_S_1_L_2_out, I0 =>  inp_feat(306), I1 =>  inp_feat(190), I2 =>  inp_feat(94), I3 =>  inp_feat(389), I4 =>  inp_feat(157), I5 =>  inp_feat(221)); 
C_30_S_1_L_3_inst : LUT6 generic map(INIT => "1000010010111100010011001110110000000000000000000000010011111010") port map( O =>C_30_S_1_L_3_out, I0 =>  inp_feat(81), I1 =>  inp_feat(153), I2 =>  inp_feat(65), I3 =>  inp_feat(224), I4 =>  inp_feat(360), I5 =>  inp_feat(84)); 
C_30_S_1_L_4_inst : LUT6 generic map(INIT => "0001000110100010101010011010001000000000001000000110000000100111") port map( O =>C_30_S_1_L_4_out, I0 =>  inp_feat(217), I1 =>  inp_feat(17), I2 =>  inp_feat(292), I3 =>  inp_feat(407), I4 =>  inp_feat(4), I5 =>  inp_feat(75)); 
C_30_S_1_L_5_inst : LUT6 generic map(INIT => "1100110101001101110011011100110000000100010001100110110000000000") port map( O =>C_30_S_1_L_5_out, I0 =>  inp_feat(269), I1 =>  inp_feat(75), I2 =>  inp_feat(162), I3 =>  inp_feat(303), I4 =>  inp_feat(130), I5 =>  inp_feat(69)); 
C_30_S_2_L_0_inst : LUT6 generic map(INIT => "0001011111011111000101110011011100010001110111111111011111111111") port map( O =>C_30_S_2_L_0_out, I0 =>  inp_feat(214), I1 =>  inp_feat(166), I2 =>  inp_feat(82), I3 =>  inp_feat(489), I4 =>  inp_feat(452), I5 =>  inp_feat(255)); 
C_30_S_2_L_1_inst : LUT6 generic map(INIT => "1100010001000011111110010111010011010000011110110111000011111000") port map( O =>C_30_S_2_L_1_out, I0 =>  inp_feat(214), I1 =>  inp_feat(361), I2 =>  inp_feat(317), I3 =>  inp_feat(278), I4 =>  inp_feat(82), I5 =>  inp_feat(360)); 
C_30_S_2_L_2_inst : LUT6 generic map(INIT => "1001100001010001000000000000000000010100001000000000000000001000") port map( O =>C_30_S_2_L_2_out, I0 =>  inp_feat(395), I1 =>  inp_feat(217), I2 =>  inp_feat(327), I3 =>  inp_feat(106), I4 =>  inp_feat(451), I5 =>  inp_feat(334)); 
C_30_S_2_L_3_inst : LUT6 generic map(INIT => "1111111100011111101111110000110100101011010000010000001000000010") port map( O =>C_30_S_2_L_3_out, I0 =>  inp_feat(204), I1 =>  inp_feat(336), I2 =>  inp_feat(306), I3 =>  inp_feat(389), I4 =>  inp_feat(325), I5 =>  inp_feat(157)); 
C_30_S_2_L_4_inst : LUT6 generic map(INIT => "1011000011110010011101001111001000000001000100001000000010100110") port map( O =>C_30_S_2_L_4_out, I0 =>  inp_feat(31), I1 =>  inp_feat(132), I2 =>  inp_feat(112), I3 =>  inp_feat(198), I4 =>  inp_feat(228), I5 =>  inp_feat(292)); 
C_30_S_2_L_5_inst : LUT6 generic map(INIT => "0100000000010001011100001011001001110010011110001111101011111011") port map( O =>C_30_S_2_L_5_out, I0 =>  inp_feat(285), I1 =>  inp_feat(17), I2 =>  inp_feat(292), I3 =>  inp_feat(82), I4 =>  inp_feat(166), I5 =>  inp_feat(93)); 
C_30_S_3_L_0_inst : LUT6 generic map(INIT => "0010111111100011000010110001111101100111111110110011111101111111") port map( O =>C_30_S_3_L_0_out, I0 =>  inp_feat(307), I1 =>  inp_feat(214), I2 =>  inp_feat(360), I3 =>  inp_feat(321), I4 =>  inp_feat(452), I5 =>  inp_feat(255)); 
C_30_S_3_L_1_inst : LUT6 generic map(INIT => "1101110110100001101001000000001001110101110001000000000001001000") port map( O =>C_30_S_3_L_1_out, I0 =>  inp_feat(255), I1 =>  inp_feat(393), I2 =>  inp_feat(132), I3 =>  inp_feat(180), I4 =>  inp_feat(316), I5 =>  inp_feat(263)); 
C_30_S_3_L_2_inst : LUT6 generic map(INIT => "1011011111010111001010100100110100000001000100000000000001000000") port map( O =>C_30_S_3_L_2_out, I0 =>  inp_feat(166), I1 =>  inp_feat(210), I2 =>  inp_feat(276), I3 =>  inp_feat(235), I4 =>  inp_feat(253), I5 =>  inp_feat(38)); 
C_30_S_3_L_3_inst : LUT6 generic map(INIT => "0010000011100011000010011111000110000000111010101111001011110001") port map( O =>C_30_S_3_L_3_out, I0 =>  inp_feat(76), I1 =>  inp_feat(278), I2 =>  inp_feat(112), I3 =>  inp_feat(93), I4 =>  inp_feat(166), I5 =>  inp_feat(82)); 
C_30_S_3_L_4_inst : LUT6 generic map(INIT => "1001011100010111110101110011000111111011000100110000000000000000") port map( O =>C_30_S_3_L_4_out, I0 =>  inp_feat(245), I1 =>  inp_feat(210), I2 =>  inp_feat(378), I3 =>  inp_feat(195), I4 =>  inp_feat(473), I5 =>  inp_feat(505)); 
C_30_S_3_L_5_inst : LUT6 generic map(INIT => "0000110010101000000000001100010011111000101100000000000000000000") port map( O =>C_30_S_3_L_5_out, I0 =>  inp_feat(478), I1 =>  inp_feat(59), I2 =>  inp_feat(81), I3 =>  inp_feat(106), I4 =>  inp_feat(473), I5 =>  inp_feat(505)); 
C_30_S_4_L_0_inst : LUT6 generic map(INIT => "1011011111110111011010100100110100000001100100000000000001000000") port map( O =>C_30_S_4_L_0_out, I0 =>  inp_feat(166), I1 =>  inp_feat(210), I2 =>  inp_feat(276), I3 =>  inp_feat(235), I4 =>  inp_feat(253), I5 =>  inp_feat(38)); 
C_30_S_4_L_1_inst : LUT6 generic map(INIT => "0000000000001101100011001100100000001010111111000000111010001100") port map( O =>C_30_S_4_L_1_out, I0 =>  inp_feat(170), I1 =>  inp_feat(317), I2 =>  inp_feat(500), I3 =>  inp_feat(82), I4 =>  inp_feat(255), I5 =>  inp_feat(367)); 
C_30_S_4_L_2_inst : LUT6 generic map(INIT => "1110001111101100110011101100100000000100000000000000100100000000") port map( O =>C_30_S_4_L_2_out, I0 =>  inp_feat(195), I1 =>  inp_feat(158), I2 =>  inp_feat(476), I3 =>  inp_feat(303), I4 =>  inp_feat(130), I5 =>  inp_feat(447)); 
C_30_S_4_L_3_inst : LUT6 generic map(INIT => "1000101011010000001010101011010000001000000010001101000110110000") port map( O =>C_30_S_4_L_3_out, I0 =>  inp_feat(346), I1 =>  inp_feat(494), I2 =>  inp_feat(88), I3 =>  inp_feat(198), I4 =>  inp_feat(228), I5 =>  inp_feat(292)); 
C_30_S_4_L_4_inst : LUT6 generic map(INIT => "0000000100010011101100010111011111010111000111110001101111110111") port map( O =>C_30_S_4_L_4_out, I0 =>  inp_feat(166), I1 =>  inp_feat(17), I2 =>  inp_feat(407), I3 =>  inp_feat(321), I4 =>  inp_feat(452), I5 =>  inp_feat(269)); 
C_30_S_4_L_5_inst : LUT6 generic map(INIT => "0100110110110101010001001011011111101000101000000000000000000000") port map( O =>C_30_S_4_L_5_out, I0 =>  inp_feat(108), I1 =>  inp_feat(86), I2 =>  inp_feat(24), I3 =>  inp_feat(189), I4 =>  inp_feat(295), I5 =>  inp_feat(400)); 
C_30_S_5_L_0_inst : LUT6 generic map(INIT => "0101000011010100001010001100101011111100011101100000000011010100") port map( O =>C_30_S_5_L_0_out, I0 =>  inp_feat(93), I1 =>  inp_feat(221), I2 =>  inp_feat(429), I3 =>  inp_feat(306), I4 =>  inp_feat(389), I5 =>  inp_feat(228)); 
C_30_S_5_L_1_inst : LUT6 generic map(INIT => "1101110100101000101100110000000000000010000001001111101000000000") port map( O =>C_30_S_5_L_1_out, I0 =>  inp_feat(470), I1 =>  inp_feat(369), I2 =>  inp_feat(357), I3 =>  inp_feat(329), I4 =>  inp_feat(508), I5 =>  inp_feat(250)); 
C_30_S_5_L_2_inst : LUT6 generic map(INIT => "0010000000001000000100000001001111111010001110001111000101110000") port map( O =>C_30_S_5_L_2_out, I0 =>  inp_feat(81), I1 =>  inp_feat(378), I2 =>  inp_feat(317), I3 =>  inp_feat(368), I4 =>  inp_feat(4), I5 =>  inp_feat(177)); 
C_30_S_5_L_3_inst : LUT6 generic map(INIT => "1010001000100000110100001001000010011100001000011001110011101100") port map( O =>C_30_S_5_L_3_out, I0 =>  inp_feat(301), I1 =>  inp_feat(70), I2 =>  inp_feat(462), I3 =>  inp_feat(24), I4 =>  inp_feat(277), I5 =>  inp_feat(8)); 
C_30_S_5_L_4_inst : LUT6 generic map(INIT => "0001010100110011110011001000000000010010000100011100010000000000") port map( O =>C_30_S_5_L_4_out, I0 =>  inp_feat(395), I1 =>  inp_feat(189), I2 =>  inp_feat(283), I3 =>  inp_feat(226), I4 =>  inp_feat(130), I5 =>  inp_feat(492)); 
C_30_S_5_L_5_inst : LUT6 generic map(INIT => "1111001101001001111100110111111000010001000000011111011100001111") port map( O =>C_30_S_5_L_5_out, I0 =>  inp_feat(229), I1 =>  inp_feat(187), I2 =>  inp_feat(446), I3 =>  inp_feat(472), I4 =>  inp_feat(437), I5 =>  inp_feat(283)); 
C_31_S_0_L_0_inst : LUT6 generic map(INIT => "0000000100000001000001010011111100010101000011110001011111111111") port map( O =>C_31_S_0_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(500), I2 =>  inp_feat(307), I3 =>  inp_feat(324), I4 =>  inp_feat(245), I5 =>  inp_feat(424)); 
C_31_S_0_L_1_inst : LUT6 generic map(INIT => "0001010100110111101111110111111110100111011111110001111111111111") port map( O =>C_31_S_0_L_1_out, I0 =>  inp_feat(46), I1 =>  inp_feat(378), I2 =>  inp_feat(17), I3 =>  inp_feat(166), I4 =>  inp_feat(280), I5 =>  inp_feat(403)); 
C_31_S_0_L_2_inst : LUT6 generic map(INIT => "0000000101101110100111111110111111111111000001010111011100010001") port map( O =>C_31_S_0_L_2_out, I0 =>  inp_feat(294), I1 =>  inp_feat(51), I2 =>  inp_feat(296), I3 =>  inp_feat(93), I4 =>  inp_feat(224), I5 =>  inp_feat(472)); 
C_31_S_0_L_3_inst : LUT6 generic map(INIT => "1010111111001011001011110000001000000001100010000000001000000000") port map( O =>C_31_S_0_L_3_out, I0 =>  inp_feat(267), I1 =>  inp_feat(17), I2 =>  inp_feat(321), I3 =>  inp_feat(170), I4 =>  inp_feat(372), I5 =>  inp_feat(413)); 
C_31_S_0_L_4_inst : LUT6 generic map(INIT => "1100010010000000000000001111001010110000111100010111000111111111") port map( O =>C_31_S_0_L_4_out, I0 =>  inp_feat(278), I1 =>  inp_feat(214), I2 =>  inp_feat(292), I3 =>  inp_feat(363), I4 =>  inp_feat(468), I5 =>  inp_feat(4)); 
C_31_S_0_L_5_inst : LUT6 generic map(INIT => "0011000100010000001101101000000011111001001100001010000010000000") port map( O =>C_31_S_0_L_5_out, I0 =>  inp_feat(47), I1 =>  inp_feat(220), I2 =>  inp_feat(180), I3 =>  inp_feat(196), I4 =>  inp_feat(468), I5 =>  inp_feat(4)); 
C_31_S_1_L_0_inst : LUT6 generic map(INIT => "0001010100110111101111110111111110100111011111110001111111111111") port map( O =>C_31_S_1_L_0_out, I0 =>  inp_feat(46), I1 =>  inp_feat(378), I2 =>  inp_feat(17), I3 =>  inp_feat(166), I4 =>  inp_feat(280), I5 =>  inp_feat(403)); 
C_31_S_1_L_1_inst : LUT6 generic map(INIT => "0000000101101110100111111110111111111111000001010111011100010001") port map( O =>C_31_S_1_L_1_out, I0 =>  inp_feat(294), I1 =>  inp_feat(51), I2 =>  inp_feat(296), I3 =>  inp_feat(93), I4 =>  inp_feat(224), I5 =>  inp_feat(472)); 
C_31_S_1_L_2_inst : LUT6 generic map(INIT => "1010111111001011001011110000001000000001100010000000001000000000") port map( O =>C_31_S_1_L_2_out, I0 =>  inp_feat(267), I1 =>  inp_feat(17), I2 =>  inp_feat(321), I3 =>  inp_feat(170), I4 =>  inp_feat(372), I5 =>  inp_feat(413)); 
C_31_S_1_L_3_inst : LUT6 generic map(INIT => "1100010010000000000000001111001010110000111100010111000111111111") port map( O =>C_31_S_1_L_3_out, I0 =>  inp_feat(278), I1 =>  inp_feat(214), I2 =>  inp_feat(292), I3 =>  inp_feat(363), I4 =>  inp_feat(468), I5 =>  inp_feat(4)); 
C_31_S_1_L_4_inst : LUT6 generic map(INIT => "0011000100010000001101101000000011111001001100001010000010000000") port map( O =>C_31_S_1_L_4_out, I0 =>  inp_feat(47), I1 =>  inp_feat(220), I2 =>  inp_feat(180), I3 =>  inp_feat(196), I4 =>  inp_feat(468), I5 =>  inp_feat(4)); 
C_31_S_1_L_5_inst : LUT6 generic map(INIT => "1001101100011111011101011111011110011001010111110000000000110111") port map( O =>C_31_S_1_L_5_out, I0 =>  inp_feat(166), I1 =>  inp_feat(360), I2 =>  inp_feat(168), I3 =>  inp_feat(424), I4 =>  inp_feat(481), I5 =>  inp_feat(63)); 
C_31_S_2_L_0_inst : LUT6 generic map(INIT => "0001000001010000011111010100001011110111000000001111011100000101") port map( O =>C_31_S_2_L_0_out, I0 =>  inp_feat(166), I1 =>  inp_feat(46), I2 =>  inp_feat(452), I3 =>  inp_feat(399), I4 =>  inp_feat(17), I5 =>  inp_feat(321)); 
C_31_S_2_L_1_inst : LUT6 generic map(INIT => "1010100001110100101011000000000010011000000000101100100011000000") port map( O =>C_31_S_2_L_1_out, I0 =>  inp_feat(110), I1 =>  inp_feat(351), I2 =>  inp_feat(399), I3 =>  inp_feat(196), I4 =>  inp_feat(82), I5 =>  inp_feat(360)); 
C_31_S_2_L_2_inst : LUT6 generic map(INIT => "0100011000100101000000100010000000111111010011111010110000000100") port map( O =>C_31_S_2_L_2_out, I0 =>  inp_feat(55), I1 =>  inp_feat(106), I2 =>  inp_feat(419), I3 =>  inp_feat(256), I4 =>  inp_feat(279), I5 =>  inp_feat(220)); 
C_31_S_2_L_3_inst : LUT6 generic map(INIT => "1101110101001010000110001100101000000001000000000000000000001000") port map( O =>C_31_S_2_L_3_out, I0 =>  inp_feat(261), I1 =>  inp_feat(39), I2 =>  inp_feat(46), I3 =>  inp_feat(177), I4 =>  inp_feat(387), I5 =>  inp_feat(432)); 
C_31_S_2_L_4_inst : LUT6 generic map(INIT => "0101010100100000011101110000001000110111101000100011111100001010") port map( O =>C_31_S_2_L_4_out, I0 =>  inp_feat(70), I1 =>  inp_feat(214), I2 =>  inp_feat(245), I3 =>  inp_feat(432), I4 =>  inp_feat(166), I5 =>  inp_feat(82)); 
C_31_S_2_L_5_inst : LUT6 generic map(INIT => "1110110011100100000110000000100000001100000000001000110010001100") port map( O =>C_31_S_2_L_5_out, I0 =>  inp_feat(135), I1 =>  inp_feat(221), I2 =>  inp_feat(130), I3 =>  inp_feat(391), I4 =>  inp_feat(121), I5 =>  inp_feat(411)); 
C_31_S_3_L_0_inst : LUT6 generic map(INIT => "0001000010100111000111011000111111000001001111110101111111111111") port map( O =>C_31_S_3_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(81), I2 =>  inp_feat(214), I3 =>  inp_feat(321), I4 =>  inp_feat(82), I5 =>  inp_feat(360)); 
C_31_S_3_L_1_inst : LUT6 generic map(INIT => "1111000000000001010101000010000000100000000101011011100001100000") port map( O =>C_31_S_3_L_1_out, I0 =>  inp_feat(423), I1 =>  inp_feat(262), I2 =>  inp_feat(454), I3 =>  inp_feat(178), I4 =>  inp_feat(321), I5 =>  inp_feat(46)); 
C_31_S_3_L_2_inst : LUT6 generic map(INIT => "0001100100010110000001110111111110010011010111110111111111111111") port map( O =>C_31_S_3_L_2_out, I0 =>  inp_feat(378), I1 =>  inp_feat(177), I2 =>  inp_feat(136), I3 =>  inp_feat(50), I4 =>  inp_feat(321), I5 =>  inp_feat(46)); 
C_31_S_3_L_3_inst : LUT6 generic map(INIT => "1000110101110001101000100000000011001101111100000000000000000000") port map( O =>C_31_S_3_L_3_out, I0 =>  inp_feat(203), I1 =>  inp_feat(180), I2 =>  inp_feat(224), I3 =>  inp_feat(173), I4 =>  inp_feat(221), I5 =>  inp_feat(411)); 
C_31_S_3_L_4_inst : LUT6 generic map(INIT => "0001000101111101010111011111111111100000000010001101000000000000") port map( O =>C_31_S_3_L_4_out, I0 =>  inp_feat(166), I1 =>  inp_feat(456), I2 =>  inp_feat(254), I3 =>  inp_feat(93), I4 =>  inp_feat(162), I5 =>  inp_feat(277)); 
C_31_S_3_L_5_inst : LUT6 generic map(INIT => "0101010100001000101010000000010011111111100011011111010001000000") port map( O =>C_31_S_3_L_5_out, I0 =>  inp_feat(21), I1 =>  inp_feat(404), I2 =>  inp_feat(114), I3 =>  inp_feat(199), I4 =>  inp_feat(481), I5 =>  inp_feat(63)); 
C_31_S_4_L_0_inst : LUT6 generic map(INIT => "1101111111011100010110010000000000001000000011000000101000000000") port map( O =>C_31_S_4_L_0_out, I0 =>  inp_feat(141), I1 =>  inp_feat(239), I2 =>  inp_feat(101), I3 =>  inp_feat(221), I4 =>  inp_feat(173), I5 =>  inp_feat(279)); 
C_31_S_4_L_1_inst : LUT6 generic map(INIT => "0001001000010010001000100000001010010000010100001101100000000000") port map( O =>C_31_S_4_L_1_out, I0 =>  inp_feat(281), I1 =>  inp_feat(94), I2 =>  inp_feat(29), I3 =>  inp_feat(454), I4 =>  inp_feat(321), I5 =>  inp_feat(46)); 
C_31_S_4_L_2_inst : LUT6 generic map(INIT => "0111101100010010010110001101011111110110000100001000100100110000") port map( O =>C_31_S_4_L_2_out, I0 =>  inp_feat(162), I1 =>  inp_feat(93), I2 =>  inp_feat(441), I3 =>  inp_feat(482), I4 =>  inp_feat(99), I5 =>  inp_feat(501)); 
C_31_S_4_L_3_inst : LUT6 generic map(INIT => "1011101100001000001111010000010010110101111101010000001000110100") port map( O =>C_31_S_4_L_3_out, I0 =>  inp_feat(120), I1 =>  inp_feat(73), I2 =>  inp_feat(63), I3 =>  inp_feat(196), I4 =>  inp_feat(434), I5 =>  inp_feat(49)); 
C_31_S_4_L_4_inst : LUT6 generic map(INIT => "0000011101001111110000100000001001100000011000000110000000000000") port map( O =>C_31_S_4_L_4_out, I0 =>  inp_feat(208), I1 =>  inp_feat(468), I2 =>  inp_feat(166), I3 =>  inp_feat(50), I4 =>  inp_feat(479), I5 =>  inp_feat(158)); 
C_31_S_4_L_5_inst : LUT6 generic map(INIT => "0100111101010101000011000111000111101000100100000000000000001000") port map( O =>C_31_S_4_L_5_out, I0 =>  inp_feat(214), I1 =>  inp_feat(307), I2 =>  inp_feat(501), I3 =>  inp_feat(166), I4 =>  inp_feat(96), I5 =>  inp_feat(40)); 
C_31_S_5_L_0_inst : LUT6 generic map(INIT => "1000011110110010100000010000000000101110111100000000000000000000") port map( O =>C_31_S_5_L_0_out, I0 =>  inp_feat(180), I1 =>  inp_feat(114), I2 =>  inp_feat(148), I3 =>  inp_feat(248), I4 =>  inp_feat(221), I5 =>  inp_feat(411)); 
C_31_S_5_L_1_inst : LUT6 generic map(INIT => "0001111000100001100100100101000010010000001111010000000111110000") port map( O =>C_31_S_5_L_1_out, I0 =>  inp_feat(394), I1 =>  inp_feat(49), I2 =>  inp_feat(448), I3 =>  inp_feat(347), I4 =>  inp_feat(0), I5 =>  inp_feat(220)); 
C_31_S_5_L_2_inst : LUT6 generic map(INIT => "0101101101000101000000001000100010111001111100111010100000001000") port map( O =>C_31_S_5_L_2_out, I0 =>  inp_feat(424), I1 =>  inp_feat(132), I2 =>  inp_feat(90), I3 =>  inp_feat(181), I4 =>  inp_feat(440), I5 =>  inp_feat(467)); 
C_31_S_5_L_3_inst : LUT6 generic map(INIT => "0100000001011000000100001111011010101000001110000000000001110000") port map( O =>C_31_S_5_L_3_out, I0 =>  inp_feat(210), I1 =>  inp_feat(119), I2 =>  inp_feat(40), I3 =>  inp_feat(321), I4 =>  inp_feat(50), I5 =>  inp_feat(275)); 
C_31_S_5_L_4_inst : LUT6 generic map(INIT => "1011111001110001000000001110001111101111011100010000000000000000") port map( O =>C_31_S_5_L_4_out, I0 =>  inp_feat(442), I1 =>  inp_feat(435), I2 =>  inp_feat(130), I3 =>  inp_feat(399), I4 =>  inp_feat(221), I5 =>  inp_feat(411)); 
C_31_S_5_L_5_inst : LUT6 generic map(INIT => "0010100000100000000110010000000111000001000000000011000101111011") port map( O =>C_31_S_5_L_5_out, I0 =>  inp_feat(282), I1 =>  inp_feat(349), I2 =>  inp_feat(162), I3 =>  inp_feat(426), I4 =>  inp_feat(89), I5 =>  inp_feat(235)); 
C_32_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000110001011100000001000001110001011101111111") port map( O =>C_32_S_0_L_0_out, I0 =>  inp_feat(378), I1 =>  inp_feat(214), I2 =>  inp_feat(307), I3 =>  inp_feat(166), I4 =>  inp_feat(245), I5 =>  inp_feat(424)); 
C_32_S_0_L_1_inst : LUT6 generic map(INIT => "0000000110000000000101011100000110000101110000011101011111000101") port map( O =>C_32_S_0_L_1_out, I0 =>  inp_feat(250), I1 =>  inp_feat(187), I2 =>  inp_feat(392), I3 =>  inp_feat(500), I4 =>  inp_feat(403), I5 =>  inp_feat(489)); 
C_32_S_0_L_2_inst : LUT6 generic map(INIT => "0010010001111111101001000000100000100000000000011010100010000000") port map( O =>C_32_S_0_L_2_out, I0 =>  inp_feat(279), I1 =>  inp_feat(31), I2 =>  inp_feat(391), I3 =>  inp_feat(226), I4 =>  inp_feat(321), I5 =>  inp_feat(360)); 
C_32_S_0_L_3_inst : LUT6 generic map(INIT => "1101100101001000110000000000000000001010000000001100000100000000") port map( O =>C_32_S_0_L_3_out, I0 =>  inp_feat(467), I1 =>  inp_feat(345), I2 =>  inp_feat(174), I3 =>  inp_feat(183), I4 =>  inp_feat(318), I5 =>  inp_feat(84)); 
C_32_S_0_L_4_inst : LUT6 generic map(INIT => "0000001000101011011000110101111100000000000000010000001100010101") port map( O =>C_32_S_0_L_4_out, I0 =>  inp_feat(245), I1 =>  inp_feat(214), I2 =>  inp_feat(166), I3 =>  inp_feat(17), I4 =>  inp_feat(321), I5 =>  inp_feat(69)); 
C_32_S_0_L_5_inst : LUT6 generic map(INIT => "1011000110010011000000000000101000000000000000000000000000000000") port map( O =>C_32_S_0_L_5_out, I0 =>  inp_feat(191), I1 =>  inp_feat(491), I2 =>  inp_feat(351), I3 =>  inp_feat(38), I4 =>  inp_feat(275), I5 =>  inp_feat(69)); 
C_32_S_1_L_0_inst : LUT6 generic map(INIT => "0000000110000000000101011100000110000101110000011101011111000101") port map( O =>C_32_S_1_L_0_out, I0 =>  inp_feat(250), I1 =>  inp_feat(187), I2 =>  inp_feat(392), I3 =>  inp_feat(500), I4 =>  inp_feat(403), I5 =>  inp_feat(489)); 
C_32_S_1_L_1_inst : LUT6 generic map(INIT => "0010010001111111101001000000100000100000000000011010100010000000") port map( O =>C_32_S_1_L_1_out, I0 =>  inp_feat(279), I1 =>  inp_feat(31), I2 =>  inp_feat(391), I3 =>  inp_feat(226), I4 =>  inp_feat(321), I5 =>  inp_feat(360)); 
C_32_S_1_L_2_inst : LUT6 generic map(INIT => "1101100101001000110000000000000000001010000000001100000100000000") port map( O =>C_32_S_1_L_2_out, I0 =>  inp_feat(467), I1 =>  inp_feat(345), I2 =>  inp_feat(174), I3 =>  inp_feat(183), I4 =>  inp_feat(318), I5 =>  inp_feat(84)); 
C_32_S_1_L_3_inst : LUT6 generic map(INIT => "0000001000101011011000110101111100000000000000010000001100010101") port map( O =>C_32_S_1_L_3_out, I0 =>  inp_feat(245), I1 =>  inp_feat(214), I2 =>  inp_feat(166), I3 =>  inp_feat(17), I4 =>  inp_feat(321), I5 =>  inp_feat(69)); 
C_32_S_1_L_4_inst : LUT6 generic map(INIT => "1011000110010011000000000000101000000000000000000000000000000000") port map( O =>C_32_S_1_L_4_out, I0 =>  inp_feat(191), I1 =>  inp_feat(491), I2 =>  inp_feat(351), I3 =>  inp_feat(38), I4 =>  inp_feat(275), I5 =>  inp_feat(69)); 
C_32_S_1_L_5_inst : LUT6 generic map(INIT => "0001110000001100011000000000000011001111001111000001110100000000") port map( O =>C_32_S_1_L_5_out, I0 =>  inp_feat(409), I1 =>  inp_feat(18), I2 =>  inp_feat(94), I3 =>  inp_feat(413), I4 =>  inp_feat(59), I5 =>  inp_feat(38)); 
C_32_S_2_L_0_inst : LUT6 generic map(INIT => "0011000111110011000000100000000011010000110101000000000011000000") port map( O =>C_32_S_2_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(383), I2 =>  inp_feat(328), I3 =>  inp_feat(324), I4 =>  inp_feat(380), I5 =>  inp_feat(360)); 
C_32_S_2_L_1_inst : LUT6 generic map(INIT => "0111000111100010100100010000000100000000000000000000000010010000") port map( O =>C_32_S_2_L_1_out, I0 =>  inp_feat(196), I1 =>  inp_feat(491), I2 =>  inp_feat(359), I3 =>  inp_feat(351), I4 =>  inp_feat(38), I5 =>  inp_feat(275)); 
C_32_S_2_L_2_inst : LUT6 generic map(INIT => "1101011111010111111001001100111100000001000000010000000100101111") port map( O =>C_32_S_2_L_2_out, I0 =>  inp_feat(500), I1 =>  inp_feat(424), I2 =>  inp_feat(17), I3 =>  inp_feat(321), I4 =>  inp_feat(255), I5 =>  inp_feat(69)); 
C_32_S_2_L_3_inst : LUT6 generic map(INIT => "0000010000000110100010100001110000000000000000000000000000100100") port map( O =>C_32_S_2_L_3_out, I0 =>  inp_feat(21), I1 =>  inp_feat(337), I2 =>  inp_feat(491), I3 =>  inp_feat(38), I4 =>  inp_feat(296), I5 =>  inp_feat(275)); 
C_32_S_2_L_4_inst : LUT6 generic map(INIT => "1110111101000000111111100000000000000000000000000011000000001000") port map( O =>C_32_S_2_L_4_out, I0 =>  inp_feat(91), I1 =>  inp_feat(120), I2 =>  inp_feat(456), I3 =>  inp_feat(183), I4 =>  inp_feat(174), I5 =>  inp_feat(348)); 
C_32_S_2_L_5_inst : LUT6 generic map(INIT => "0000010000010011000010000110000100000000000000000000000001000000") port map( O =>C_32_S_2_L_5_out, I0 =>  inp_feat(96), I1 =>  inp_feat(359), I2 =>  inp_feat(142), I3 =>  inp_feat(408), I4 =>  inp_feat(351), I5 =>  inp_feat(275)); 
C_32_S_3_L_0_inst : LUT6 generic map(INIT => "1000000101010010010100010000100100000000000000000000000000001100") port map( O =>C_32_S_3_L_0_out, I0 =>  inp_feat(491), I1 =>  inp_feat(359), I2 =>  inp_feat(408), I3 =>  inp_feat(96), I4 =>  inp_feat(38), I5 =>  inp_feat(275)); 
C_32_S_3_L_1_inst : LUT6 generic map(INIT => "0000001101110110101100100010001000000001000001100000001011000000") port map( O =>C_32_S_3_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(321), I2 =>  inp_feat(300), I3 =>  inp_feat(22), I4 =>  inp_feat(184), I5 =>  inp_feat(380)); 
C_32_S_3_L_2_inst : LUT6 generic map(INIT => "1101001011000000100000000000000000000000000001000000000011000000") port map( O =>C_32_S_3_L_2_out, I0 =>  inp_feat(376), I1 =>  inp_feat(201), I2 =>  inp_feat(349), I3 =>  inp_feat(362), I4 =>  inp_feat(184), I5 =>  inp_feat(380)); 
C_32_S_3_L_3_inst : LUT6 generic map(INIT => "0001000101001011101111110111111100000000000100010000000100010111") port map( O =>C_32_S_3_L_3_out, I0 =>  inp_feat(324), I1 =>  inp_feat(278), I2 =>  inp_feat(210), I3 =>  inp_feat(468), I4 =>  inp_feat(4), I5 =>  inp_feat(69)); 
C_32_S_3_L_4_inst : LUT6 generic map(INIT => "1000000100001001100000001000110000000000000010000000100010001000") port map( O =>C_32_S_3_L_4_out, I0 =>  inp_feat(488), I1 =>  inp_feat(312), I2 =>  inp_feat(17), I3 =>  inp_feat(166), I4 =>  inp_feat(132), I5 =>  inp_feat(69)); 
C_32_S_3_L_5_inst : LUT6 generic map(INIT => "0100000001010100000010001111000000000000000000000001000000000100") port map( O =>C_32_S_3_L_5_out, I0 =>  inp_feat(408), I1 =>  inp_feat(335), I2 =>  inp_feat(7), I3 =>  inp_feat(491), I4 =>  inp_feat(296), I5 =>  inp_feat(275)); 
C_32_S_4_L_0_inst : LUT6 generic map(INIT => "0011010100000101000101110000001101010111000000011111111100100011") port map( O =>C_32_S_4_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(82), I2 =>  inp_feat(46), I3 =>  inp_feat(2), I4 =>  inp_feat(280), I5 =>  inp_feat(406)); 
C_32_S_4_L_1_inst : LUT6 generic map(INIT => "1101110111001100010000100000110000000000000001000000000011000000") port map( O =>C_32_S_4_L_1_out, I0 =>  inp_feat(126), I1 =>  inp_feat(76), I2 =>  inp_feat(120), I3 =>  inp_feat(441), I4 =>  inp_feat(109), I5 =>  inp_feat(348)); 
C_32_S_4_L_2_inst : LUT6 generic map(INIT => "0001001010010000001100001101000000000000000000000001000000001000") port map( O =>C_32_S_4_L_2_out, I0 =>  inp_feat(82), I1 =>  inp_feat(50), I2 =>  inp_feat(158), I3 =>  inp_feat(491), I4 =>  inp_feat(296), I5 =>  inp_feat(275)); 
C_32_S_4_L_3_inst : LUT6 generic map(INIT => "1111001011110000010100000011000000010000000000001000000000000000") port map( O =>C_32_S_4_L_3_out, I0 =>  inp_feat(406), I1 =>  inp_feat(166), I2 =>  inp_feat(317), I3 =>  inp_feat(322), I4 =>  inp_feat(33), I5 =>  inp_feat(59)); 
C_32_S_4_L_4_inst : LUT6 generic map(INIT => "0000100001000010000100011011000000000000000000000001000000001000") port map( O =>C_32_S_4_L_4_out, I0 =>  inp_feat(501), I1 =>  inp_feat(392), I2 =>  inp_feat(153), I3 =>  inp_feat(389), I4 =>  inp_feat(38), I5 =>  inp_feat(275)); 
C_32_S_4_L_5_inst : LUT6 generic map(INIT => "1000110011010000100100001011000100000000000000000000001000000000") port map( O =>C_32_S_4_L_5_out, I0 =>  inp_feat(176), I1 =>  inp_feat(189), I2 =>  inp_feat(38), I3 =>  inp_feat(142), I4 =>  inp_feat(296), I5 =>  inp_feat(275)); 
C_32_S_5_L_0_inst : LUT6 generic map(INIT => "0110111110000000000000101111000101010101001000000000000011000001") port map( O =>C_32_S_5_L_0_out, I0 =>  inp_feat(177), I1 =>  inp_feat(307), I2 =>  inp_feat(162), I3 =>  inp_feat(215), I4 =>  inp_feat(187), I5 =>  inp_feat(1)); 
C_32_S_5_L_1_inst : LUT6 generic map(INIT => "0000110010010110000000001011110000001010000001000000000010000110") port map( O =>C_32_S_5_L_1_out, I0 =>  inp_feat(141), I1 =>  inp_feat(467), I2 =>  inp_feat(164), I3 =>  inp_feat(194), I4 =>  inp_feat(94), I5 =>  inp_feat(417)); 
C_32_S_5_L_2_inst : LUT6 generic map(INIT => "0001000000000001111101110000001111010111000000001111111100010011") port map( O =>C_32_S_5_L_2_out, I0 =>  inp_feat(458), I1 =>  inp_feat(166), I2 =>  inp_feat(424), I3 =>  inp_feat(270), I4 =>  inp_feat(210), I5 =>  inp_feat(70)); 
C_32_S_5_L_3_inst : LUT6 generic map(INIT => "1111110000101111010000000100110000010000011000011001001000000000") port map( O =>C_32_S_5_L_3_out, I0 =>  inp_feat(242), I1 =>  inp_feat(113), I2 =>  inp_feat(101), I3 =>  inp_feat(187), I4 =>  inp_feat(133), I5 =>  inp_feat(83)); 
C_32_S_5_L_4_inst : LUT6 generic map(INIT => "0000000000101110000000000010101100000000000000110000001000101011") port map( O =>C_32_S_5_L_4_out, I0 =>  inp_feat(292), I1 =>  inp_feat(278), I2 =>  inp_feat(17), I3 =>  inp_feat(166), I4 =>  inp_feat(132), I5 =>  inp_feat(69)); 
C_32_S_5_L_5_inst : LUT6 generic map(INIT => "1101111011011001000100011111011100000000000100000001010110010001") port map( O =>C_32_S_5_L_5_out, I0 =>  inp_feat(17), I1 =>  inp_feat(177), I2 =>  inp_feat(122), I3 =>  inp_feat(130), I4 =>  inp_feat(424), I5 =>  inp_feat(366)); 
C_33_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000010111011100000001000101110000011111111111") port map( O =>C_33_S_0_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(214), I2 =>  inp_feat(166), I3 =>  inp_feat(307), I4 =>  inp_feat(17), I5 =>  inp_feat(321)); 
C_33_S_0_L_1_inst : LUT6 generic map(INIT => "0000000100001111100000010001111110000000100011111111001101111111") port map( O =>C_33_S_0_L_1_out, I0 =>  inp_feat(44), I1 =>  inp_feat(182), I2 =>  inp_feat(211), I3 =>  inp_feat(239), I4 =>  inp_feat(403), I5 =>  inp_feat(489)); 
C_33_S_0_L_2_inst : LUT6 generic map(INIT => "1101010100000011111101110100000000000010000000100100000001000000") port map( O =>C_33_S_0_L_2_out, I0 =>  inp_feat(46), I1 =>  inp_feat(280), I2 =>  inp_feat(257), I3 =>  inp_feat(432), I4 =>  inp_feat(418), I5 =>  inp_feat(183)); 
C_33_S_0_L_3_inst : LUT6 generic map(INIT => "0000000100110010110101110000000010010001110010001111111100000000") port map( O =>C_33_S_0_L_3_out, I0 =>  inp_feat(166), I1 =>  inp_feat(321), I2 =>  inp_feat(70), I3 =>  inp_feat(197), I4 =>  inp_feat(407), I5 =>  inp_feat(463)); 
C_33_S_0_L_4_inst : LUT6 generic map(INIT => "1100010100011111111101110101111100010111100111110001111101111111") port map( O =>C_33_S_0_L_4_out, I0 =>  inp_feat(46), I1 =>  inp_feat(162), I2 =>  inp_feat(324), I3 =>  inp_feat(177), I4 =>  inp_feat(321), I5 =>  inp_feat(138)); 
C_33_S_0_L_5_inst : LUT6 generic map(INIT => "1111101011000101000100001111001100010000110100000000000000000000") port map( O =>C_33_S_0_L_5_out, I0 =>  inp_feat(227), I1 =>  inp_feat(249), I2 =>  inp_feat(147), I3 =>  inp_feat(78), I4 =>  inp_feat(312), I5 =>  inp_feat(418)); 
C_33_S_1_L_0_inst : LUT6 generic map(INIT => "0000000100001111000000100011111111000000010011111010001101111111") port map( O =>C_33_S_1_L_0_out, I0 =>  inp_feat(303), I1 =>  inp_feat(182), I2 =>  inp_feat(211), I3 =>  inp_feat(239), I4 =>  inp_feat(403), I5 =>  inp_feat(489)); 
C_33_S_1_L_1_inst : LUT6 generic map(INIT => "1100111001000010001010100000101100000100110000000000000000000010") port map( O =>C_33_S_1_L_1_out, I0 =>  inp_feat(334), I1 =>  inp_feat(424), I2 =>  inp_feat(245), I3 =>  inp_feat(248), I4 =>  inp_feat(257), I5 =>  inp_feat(183)); 
C_33_S_1_L_2_inst : LUT6 generic map(INIT => "1011000000000000010111111000100000001000000000000000011011110000") port map( O =>C_33_S_1_L_2_out, I0 =>  inp_feat(405), I1 =>  inp_feat(106), I2 =>  inp_feat(313), I3 =>  inp_feat(20), I4 =>  inp_feat(78), I5 =>  inp_feat(52)); 
C_33_S_1_L_3_inst : LUT6 generic map(INIT => "1100000100111111000000001001011000000011000100010000000000000000") port map( O =>C_33_S_1_L_3_out, I0 =>  inp_feat(245), I1 =>  inp_feat(307), I2 =>  inp_feat(166), I3 =>  inp_feat(257), I4 =>  inp_feat(112), I5 =>  inp_feat(418)); 
C_33_S_1_L_4_inst : LUT6 generic map(INIT => "0001000011010001011100111111011100010010010100011111001111111111") port map( O =>C_33_S_1_L_4_out, I0 =>  inp_feat(338), I1 =>  inp_feat(177), I2 =>  inp_feat(306), I3 =>  inp_feat(307), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_1_L_5_inst : LUT6 generic map(INIT => "1111111110110110001101111010000000000100000000010000000000000000") port map( O =>C_33_S_1_L_5_out, I0 =>  inp_feat(279), I1 =>  inp_feat(30), I2 =>  inp_feat(419), I3 =>  inp_feat(424), I4 =>  inp_feat(70), I5 =>  inp_feat(234)); 
C_33_S_2_L_0_inst : LUT6 generic map(INIT => "0000000010010111001000110111111111110010000101110000111111111111") port map( O =>C_33_S_2_L_0_out, I0 =>  inp_feat(360), I1 =>  inp_feat(378), I2 =>  inp_feat(46), I3 =>  inp_feat(245), I4 =>  inp_feat(324), I5 =>  inp_feat(403)); 
C_33_S_2_L_1_inst : LUT6 generic map(INIT => "0111111100010111001100100000000000100011000000011011001000000000") port map( O =>C_33_S_2_L_1_out, I0 =>  inp_feat(394), I1 =>  inp_feat(100), I2 =>  inp_feat(440), I3 =>  inp_feat(14), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_2_L_2_inst : LUT6 generic map(INIT => "0010001100010111111000100000001110011101010001111000110011000000") port map( O =>C_33_S_2_L_2_out, I0 =>  inp_feat(70), I1 =>  inp_feat(324), I2 =>  inp_feat(307), I3 =>  inp_feat(500), I4 =>  inp_feat(111), I5 =>  inp_feat(471)); 
C_33_S_2_L_3_inst : LUT6 generic map(INIT => "1101111110000101010111110010000101010101010101010000011000011000") port map( O =>C_33_S_2_L_3_out, I0 =>  inp_feat(307), I1 =>  inp_feat(404), I2 =>  inp_feat(361), I3 =>  inp_feat(173), I4 =>  inp_feat(273), I5 =>  inp_feat(65)); 
C_33_S_2_L_4_inst : LUT6 generic map(INIT => "1011000100010011001110010000000000000000000000000000000000000001") port map( O =>C_33_S_2_L_4_out, I0 =>  inp_feat(353), I1 =>  inp_feat(44), I2 =>  inp_feat(470), I3 =>  inp_feat(173), I4 =>  inp_feat(13), I5 =>  inp_feat(112)); 
C_33_S_2_L_5_inst : LUT6 generic map(INIT => "0000100100101010000000100000101110010010111010100011101010101111") port map( O =>C_33_S_2_L_5_out, I0 =>  inp_feat(426), I1 =>  inp_feat(224), I2 =>  inp_feat(458), I3 =>  inp_feat(166), I4 =>  inp_feat(17), I5 =>  inp_feat(321)); 
C_33_S_3_L_0_inst : LUT6 generic map(INIT => "0111011100010111001100110000000000100011000000011011001000000000") port map( O =>C_33_S_3_L_0_out, I0 =>  inp_feat(394), I1 =>  inp_feat(100), I2 =>  inp_feat(440), I3 =>  inp_feat(14), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_3_L_1_inst : LUT6 generic map(INIT => "1100010101100111110000010000111100000001001011110001011101111111") port map( O =>C_33_S_3_L_1_out, I0 =>  inp_feat(468), I1 =>  inp_feat(210), I2 =>  inp_feat(245), I3 =>  inp_feat(324), I4 =>  inp_feat(162), I5 =>  inp_feat(424)); 
C_33_S_3_L_2_inst : LUT6 generic map(INIT => "0100011110000111001101110101111100000011001111110011011111111111") port map( O =>C_33_S_3_L_2_out, I0 =>  inp_feat(321), I1 =>  inp_feat(4), I2 =>  inp_feat(278), I3 =>  inp_feat(324), I4 =>  inp_feat(162), I5 =>  inp_feat(424)); 
C_33_S_3_L_3_inst : LUT6 generic map(INIT => "1000101010010000011100001101010010110000001100111111000111110111") port map( O =>C_33_S_3_L_3_out, I0 =>  inp_feat(363), I1 =>  inp_feat(4), I2 =>  inp_feat(292), I3 =>  inp_feat(46), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_3_L_4_inst : LUT6 generic map(INIT => "0000001100000011100100110011111100010001001111110001111111111111") port map( O =>C_33_S_3_L_4_out, I0 =>  inp_feat(500), I1 =>  inp_feat(82), I2 =>  inp_feat(4), I3 =>  inp_feat(324), I4 =>  inp_feat(278), I5 =>  inp_feat(424)); 
C_33_S_3_L_5_inst : LUT6 generic map(INIT => "1000100000000011000101110111111100010001011011110111111111111111") port map( O =>C_33_S_3_L_5_out, I0 =>  inp_feat(378), I1 =>  inp_feat(82), I2 =>  inp_feat(4), I3 =>  inp_feat(324), I4 =>  inp_feat(278), I5 =>  inp_feat(424)); 
C_33_S_4_L_0_inst : LUT6 generic map(INIT => "0101011000010111010101000000000010100011000010011111001000000000") port map( O =>C_33_S_4_L_0_out, I0 =>  inp_feat(386), I1 =>  inp_feat(100), I2 =>  inp_feat(440), I3 =>  inp_feat(14), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_4_L_1_inst : LUT6 generic map(INIT => "1000110011010000001111000111100000011000011100000111100001110011") port map( O =>C_33_S_4_L_1_out, I0 =>  inp_feat(378), I1 =>  inp_feat(245), I2 =>  inp_feat(116), I3 =>  inp_feat(46), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_4_L_2_inst : LUT6 generic map(INIT => "1000110110100011100000010000111100000011001011110001010101111111") port map( O =>C_33_S_4_L_2_out, I0 =>  inp_feat(500), I1 =>  inp_feat(210), I2 =>  inp_feat(245), I3 =>  inp_feat(324), I4 =>  inp_feat(162), I5 =>  inp_feat(424)); 
C_33_S_4_L_3_inst : LUT6 generic map(INIT => "0000000110000010000101111001000010010011000000000111111100011000") port map( O =>C_33_S_4_L_3_out, I0 =>  inp_feat(214), I1 =>  inp_feat(166), I2 =>  inp_feat(255), I3 =>  inp_feat(473), I4 =>  inp_feat(177), I5 =>  inp_feat(424)); 
C_33_S_4_L_4_inst : LUT6 generic map(INIT => "1010101110000011000110110011111100010001011111110001111111111111") port map( O =>C_33_S_4_L_4_out, I0 =>  inp_feat(500), I1 =>  inp_feat(82), I2 =>  inp_feat(4), I3 =>  inp_feat(324), I4 =>  inp_feat(278), I5 =>  inp_feat(424)); 
C_33_S_4_L_5_inst : LUT6 generic map(INIT => "0000001000000010100010100010101001000010001010100010101011101010") port map( O =>C_33_S_4_L_5_out, I0 =>  inp_feat(335), I1 =>  inp_feat(237), I2 =>  inp_feat(4), I3 =>  inp_feat(324), I4 =>  inp_feat(278), I5 =>  inp_feat(424)); 
C_33_S_5_L_0_inst : LUT6 generic map(INIT => "1010111000010011111101100000000010100011000010011111001000000000") port map( O =>C_33_S_5_L_0_out, I0 =>  inp_feat(386), I1 =>  inp_feat(100), I2 =>  inp_feat(440), I3 =>  inp_feat(14), I4 =>  inp_feat(360), I5 =>  inp_feat(424)); 
C_33_S_5_L_1_inst : LUT6 generic map(INIT => "0000000100000010000100111101000000010011000000000111111100011000") port map( O =>C_33_S_5_L_1_out, I0 =>  inp_feat(214), I1 =>  inp_feat(166), I2 =>  inp_feat(255), I3 =>  inp_feat(473), I4 =>  inp_feat(177), I5 =>  inp_feat(424)); 
C_33_S_5_L_2_inst : LUT6 generic map(INIT => "0101000110101101000111010010001111111110111011100101000000011110") port map( O =>C_33_S_5_L_2_out, I0 =>  inp_feat(190), I1 =>  inp_feat(47), I2 =>  inp_feat(375), I3 =>  inp_feat(78), I4 =>  inp_feat(438), I5 =>  inp_feat(483)); 
C_33_S_5_L_3_inst : LUT6 generic map(INIT => "1000000110000111001011110111111100000011101111110001011101111111") port map( O =>C_33_S_5_L_3_out, I0 =>  inp_feat(500), I1 =>  inp_feat(278), I2 =>  inp_feat(4), I3 =>  inp_feat(324), I4 =>  inp_feat(177), I5 =>  inp_feat(424)); 
C_33_S_5_L_4_inst : LUT6 generic map(INIT => "0000110111100111100000010000111100100011001011110001010101111111") port map( O =>C_33_S_5_L_4_out, I0 =>  inp_feat(500), I1 =>  inp_feat(210), I2 =>  inp_feat(245), I3 =>  inp_feat(324), I4 =>  inp_feat(162), I5 =>  inp_feat(424)); 
C_33_S_5_L_5_inst : LUT6 generic map(INIT => "1100100100010001000100010000111100010011010101110111011111111111") port map( O =>C_33_S_5_L_5_out, I0 =>  inp_feat(378), I1 =>  inp_feat(500), I2 =>  inp_feat(224), I3 =>  inp_feat(324), I4 =>  inp_feat(162), I5 =>  inp_feat(424)); 
C_34_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111100111111001100100011111110111010001110100010000000") port map( O =>C_34_S_0_L_0_out, I0 =>  inp_feat(255), I1 =>  inp_feat(214), I2 =>  inp_feat(307), I3 =>  inp_feat(166), I4 =>  inp_feat(245), I5 =>  inp_feat(424)); 
C_34_S_0_L_1_inst : LUT6 generic map(INIT => "1111110110110110111011000000001000000001000010100000110000000100") port map( O =>C_34_S_0_L_1_out, I0 =>  inp_feat(458), I1 =>  inp_feat(307), I2 =>  inp_feat(250), I3 =>  inp_feat(214), I4 =>  inp_feat(136), I5 =>  inp_feat(321)); 
C_34_S_0_L_2_inst : LUT6 generic map(INIT => "0000110111000101101111011000110011101000100010001110100010101000") port map( O =>C_34_S_0_L_2_out, I0 =>  inp_feat(360), I1 =>  inp_feat(21), I2 =>  inp_feat(30), I3 =>  inp_feat(292), I4 =>  inp_feat(98), I5 =>  inp_feat(183)); 
C_34_S_0_L_3_inst : LUT6 generic map(INIT => "1101010111011111010100000100110001010011110111110101001000001011") port map( O =>C_34_S_0_L_3_out, I0 =>  inp_feat(350), I1 =>  inp_feat(360), I2 =>  inp_feat(454), I3 =>  inp_feat(468), I4 =>  inp_feat(4), I5 =>  inp_feat(262)); 
C_34_S_0_L_4_inst : LUT6 generic map(INIT => "1100001001111001100110000001110001011011000101110001100000000000") port map( O =>C_34_S_0_L_4_out, I0 =>  inp_feat(248), I1 =>  inp_feat(190), I2 =>  inp_feat(226), I3 =>  inp_feat(321), I4 =>  inp_feat(468), I5 =>  inp_feat(82)); 
C_34_S_0_L_5_inst : LUT6 generic map(INIT => "0000101000101011011111100011001111111111001111110011111100010011") port map( O =>C_34_S_0_L_5_out, I0 =>  inp_feat(59), I1 =>  inp_feat(395), I2 =>  inp_feat(28), I3 =>  inp_feat(24), I4 =>  inp_feat(405), I5 =>  inp_feat(116)); 
C_34_S_1_L_0_inst : LUT6 generic map(INIT => "1111110110110110111011000000001000000001000010100000110000000100") port map( O =>C_34_S_1_L_0_out, I0 =>  inp_feat(458), I1 =>  inp_feat(307), I2 =>  inp_feat(250), I3 =>  inp_feat(214), I4 =>  inp_feat(136), I5 =>  inp_feat(321)); 
C_34_S_1_L_1_inst : LUT6 generic map(INIT => "0000110111000101101111011000110011101000100010001110100010101000") port map( O =>C_34_S_1_L_1_out, I0 =>  inp_feat(360), I1 =>  inp_feat(21), I2 =>  inp_feat(30), I3 =>  inp_feat(292), I4 =>  inp_feat(98), I5 =>  inp_feat(183)); 
C_34_S_1_L_2_inst : LUT6 generic map(INIT => "1101010111011111010100000100110001010011110111110101001000001011") port map( O =>C_34_S_1_L_2_out, I0 =>  inp_feat(350), I1 =>  inp_feat(360), I2 =>  inp_feat(454), I3 =>  inp_feat(468), I4 =>  inp_feat(4), I5 =>  inp_feat(262)); 
C_34_S_1_L_3_inst : LUT6 generic map(INIT => "1100001001111001100110000001110001011011000101110001100000000000") port map( O =>C_34_S_1_L_3_out, I0 =>  inp_feat(248), I1 =>  inp_feat(190), I2 =>  inp_feat(226), I3 =>  inp_feat(321), I4 =>  inp_feat(468), I5 =>  inp_feat(82)); 
C_34_S_1_L_4_inst : LUT6 generic map(INIT => "0000101000101011011111100011001111111111001111110011111100010011") port map( O =>C_34_S_1_L_4_out, I0 =>  inp_feat(59), I1 =>  inp_feat(395), I2 =>  inp_feat(28), I3 =>  inp_feat(24), I4 =>  inp_feat(405), I5 =>  inp_feat(116)); 
C_34_S_1_L_5_inst : LUT6 generic map(INIT => "1010110010001000011011101101110011111110101010001111111001001000") port map( O =>C_34_S_1_L_5_out, I0 =>  inp_feat(50), I1 =>  inp_feat(166), I2 =>  inp_feat(300), I3 =>  inp_feat(208), I4 =>  inp_feat(434), I5 =>  inp_feat(266)); 
C_34_S_2_L_0_inst : LUT6 generic map(INIT => "1111111110100011001111000000110001101100100011100000100000000000") port map( O =>C_34_S_2_L_0_out, I0 =>  inp_feat(166), I1 =>  inp_feat(300), I2 =>  inp_feat(454), I3 =>  inp_feat(4), I4 =>  inp_feat(500), I5 =>  inp_feat(82)); 
C_34_S_2_L_1_inst : LUT6 generic map(INIT => "1010000000011100111011100110011010100000111010001111101010000000") port map( O =>C_34_S_2_L_1_out, I0 =>  inp_feat(403), I1 =>  inp_feat(321), I2 =>  inp_feat(17), I3 =>  inp_feat(30), I4 =>  inp_feat(98), I5 =>  inp_feat(418)); 
C_34_S_2_L_2_inst : LUT6 generic map(INIT => "0100101000001000000111111110111011111101111000001111111111001000") port map( O =>C_34_S_2_L_2_out, I0 =>  inp_feat(265), I1 =>  inp_feat(463), I2 =>  inp_feat(276), I3 =>  inp_feat(208), I4 =>  inp_feat(434), I5 =>  inp_feat(266)); 
C_34_S_2_L_3_inst : LUT6 generic map(INIT => "1110000101001110111011000001101110101010110011101111111011110010") port map( O =>C_34_S_2_L_3_out, I0 =>  inp_feat(255), I1 =>  inp_feat(363), I2 =>  inp_feat(122), I3 =>  inp_feat(267), I4 =>  inp_feat(478), I5 =>  inp_feat(486)); 
C_34_S_2_L_4_inst : LUT6 generic map(INIT => "1011111101010111111111110101101100001010001011001100101010101000") port map( O =>C_34_S_2_L_4_out, I0 =>  inp_feat(162), I1 =>  inp_feat(290), I2 =>  inp_feat(7), I3 =>  inp_feat(24), I4 =>  inp_feat(26), I5 =>  inp_feat(324)); 
C_34_S_2_L_5_inst : LUT6 generic map(INIT => "0001111001010111111011000111101011101011111111001110100010100000") port map( O =>C_34_S_2_L_5_out, I0 =>  inp_feat(338), I1 =>  inp_feat(235), I2 =>  inp_feat(56), I3 =>  inp_feat(141), I4 =>  inp_feat(158), I5 =>  inp_feat(116)); 
C_34_S_3_L_0_inst : LUT6 generic map(INIT => "1111101110110011111100110011001111010010101000111011000100000000") port map( O =>C_34_S_3_L_0_out, I0 =>  inp_feat(361), I1 =>  inp_feat(230), I2 =>  inp_feat(50), I3 =>  inp_feat(321), I4 =>  inp_feat(360), I5 =>  inp_feat(82)); 
C_34_S_3_L_1_inst : LUT6 generic map(INIT => "0100011000101111011011110010001011111111111111000111010011110100") port map( O =>C_34_S_3_L_1_out, I0 =>  inp_feat(11), I1 =>  inp_feat(455), I2 =>  inp_feat(399), I3 =>  inp_feat(149), I4 =>  inp_feat(41), I5 =>  inp_feat(486)); 
C_34_S_3_L_2_inst : LUT6 generic map(INIT => "1101110110111101101000110011111100010010000000111011001011111111") port map( O =>C_34_S_3_L_2_out, I0 =>  inp_feat(417), I1 =>  inp_feat(127), I2 =>  inp_feat(173), I3 =>  inp_feat(373), I4 =>  inp_feat(182), I5 =>  inp_feat(403)); 
C_34_S_3_L_3_inst : LUT6 generic map(INIT => "0100000110100111000011001110101110001110011010110000110010101011") port map( O =>C_34_S_3_L_3_out, I0 =>  inp_feat(255), I1 =>  inp_feat(324), I2 =>  inp_feat(83), I3 =>  inp_feat(7), I4 =>  inp_feat(332), I5 =>  inp_feat(416)); 
C_34_S_3_L_4_inst : LUT6 generic map(INIT => "1100100011010010101010001100001001100011111010000000000011011101") port map( O =>C_34_S_3_L_4_out, I0 =>  inp_feat(50), I1 =>  inp_feat(156), I2 =>  inp_feat(267), I3 =>  inp_feat(440), I4 =>  inp_feat(245), I5 =>  inp_feat(416)); 
C_34_S_3_L_5_inst : LUT6 generic map(INIT => "0001111011111100000101111110111010111110111111001111111111111110") port map( O =>C_34_S_3_L_5_out, I0 =>  inp_feat(107), I1 =>  inp_feat(460), I2 =>  inp_feat(69), I3 =>  inp_feat(98), I4 =>  inp_feat(183), I5 =>  inp_feat(316)); 
C_34_S_4_L_0_inst : LUT6 generic map(INIT => "0011001000101011111101101011111111010101111111001111111100011111") port map( O =>C_34_S_4_L_0_out, I0 =>  inp_feat(389), I1 =>  inp_feat(508), I2 =>  inp_feat(472), I3 =>  inp_feat(144), I4 =>  inp_feat(182), I5 =>  inp_feat(422)); 
C_34_S_4_L_1_inst : LUT6 generic map(INIT => "1011001101011111111111011001001010111011111111111111111100001101") port map( O =>C_34_S_4_L_1_out, I0 =>  inp_feat(447), I1 =>  inp_feat(322), I2 =>  inp_feat(375), I3 =>  inp_feat(469), I4 =>  inp_feat(96), I5 =>  inp_feat(496)); 
C_34_S_4_L_2_inst : LUT6 generic map(INIT => "0010001011011000011100110100011011111011111110100010101110101010") port map( O =>C_34_S_4_L_2_out, I0 =>  inp_feat(171), I1 =>  inp_feat(317), I2 =>  inp_feat(162), I3 =>  inp_feat(369), I4 =>  inp_feat(269), I5 =>  inp_feat(496)); 
C_34_S_4_L_3_inst : LUT6 generic map(INIT => "1110111010100011111101101110011001010111111101110001000110000010") port map( O =>C_34_S_4_L_3_out, I0 =>  inp_feat(126), I1 =>  inp_feat(179), I2 =>  inp_feat(283), I3 =>  inp_feat(464), I4 =>  inp_feat(211), I5 =>  inp_feat(226)); 
C_34_S_4_L_4_inst : LUT6 generic map(INIT => "0011011011010010011011111111000011111010100000101110011110000000") port map( O =>C_34_S_4_L_4_out, I0 =>  inp_feat(148), I1 =>  inp_feat(316), I2 =>  inp_feat(166), I3 =>  inp_feat(416), I4 =>  inp_feat(226), I5 =>  inp_feat(38)); 
C_34_S_4_L_5_inst : LUT6 generic map(INIT => "1010001010111001001011101111100011111111111111011011000011111111") port map( O =>C_34_S_4_L_5_out, I0 =>  inp_feat(468), I1 =>  inp_feat(44), I2 =>  inp_feat(503), I3 =>  inp_feat(182), I4 =>  inp_feat(459), I5 =>  inp_feat(127)); 
C_34_S_5_L_0_inst : LUT6 generic map(INIT => "0001110010101110001010001111001111111111101010111010010011111111") port map( O =>C_34_S_5_L_0_out, I0 =>  inp_feat(156), I1 =>  inp_feat(500), I2 =>  inp_feat(46), I3 =>  inp_feat(330), I4 =>  inp_feat(195), I5 =>  inp_feat(127)); 
C_34_S_5_L_1_inst : LUT6 generic map(INIT => "1111101001101011100110101110101111111110111000001111111111111001") port map( O =>C_34_S_5_L_1_out, I0 =>  inp_feat(226), I1 =>  inp_feat(461), I2 =>  inp_feat(339), I3 =>  inp_feat(88), I4 =>  inp_feat(290), I5 =>  inp_feat(126)); 
C_34_S_5_L_2_inst : LUT6 generic map(INIT => "0011101101010001000001011101111111111111110111110001011101011111") port map( O =>C_34_S_5_L_2_out, I0 =>  inp_feat(489), I1 =>  inp_feat(170), I2 =>  inp_feat(270), I3 =>  inp_feat(391), I4 =>  inp_feat(59), I5 =>  inp_feat(241)); 
C_34_S_5_L_3_inst : LUT6 generic map(INIT => "1110111011101101111000111101001100101100110111001110110011001000") port map( O =>C_34_S_5_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(255), I2 =>  inp_feat(370), I3 =>  inp_feat(486), I4 =>  inp_feat(39), I5 =>  inp_feat(205)); 
C_34_S_5_L_4_inst : LUT6 generic map(INIT => "0100001101010101011101101111001101010010000100010111110011111111") port map( O =>C_34_S_5_L_4_out, I0 =>  inp_feat(434), I1 =>  inp_feat(386), I2 =>  inp_feat(195), I3 =>  inp_feat(372), I4 =>  inp_feat(183), I5 =>  inp_feat(152)); 
C_34_S_5_L_5_inst : LUT6 generic map(INIT => "1011101111010111011100111111111101111110111101101101111111111111") port map( O =>C_34_S_5_L_5_out, I0 =>  inp_feat(49), I1 =>  inp_feat(301), I2 =>  inp_feat(376), I3 =>  inp_feat(121), I4 =>  inp_feat(36), I5 =>  inp_feat(152)); 
C_35_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111101110111110101100100011101110111010001100000000000000") port map( O =>C_35_S_0_L_0_out, I0 =>  inp_feat(458), I1 =>  inp_feat(324), I2 =>  inp_feat(210), I3 =>  inp_feat(321), I4 =>  inp_feat(245), I5 =>  inp_feat(424)); 
C_35_S_0_L_1_inst : LUT6 generic map(INIT => "1111100110110010000000100000110000000000000000100011111000010000") port map( O =>C_35_S_0_L_1_out, I0 =>  inp_feat(493), I1 =>  inp_feat(429), I2 =>  inp_feat(226), I3 =>  inp_feat(162), I4 =>  inp_feat(280), I5 =>  inp_feat(321)); 
C_35_S_0_L_2_inst : LUT6 generic map(INIT => "1100011011111010111111101010001000000011101100001011000000000000") port map( O =>C_35_S_0_L_2_out, I0 =>  inp_feat(162), I1 =>  inp_feat(91), I2 =>  inp_feat(360), I3 =>  inp_feat(214), I4 =>  inp_feat(17), I5 =>  inp_feat(307)); 
C_35_S_0_L_3_inst : LUT6 generic map(INIT => "1011001110111000100001101111101001110110111000110000110111010100") port map( O =>C_35_S_0_L_3_out, I0 =>  inp_feat(162), I1 =>  inp_feat(235), I2 =>  inp_feat(394), I3 =>  inp_feat(264), I4 =>  inp_feat(468), I5 =>  inp_feat(4)); 
C_35_S_0_L_4_inst : LUT6 generic map(INIT => "1111100011111100011001000110010000000000000101001111010000110000") port map( O =>C_35_S_0_L_4_out, I0 =>  inp_feat(185), I1 =>  inp_feat(177), I2 =>  inp_feat(166), I3 =>  inp_feat(320), I4 =>  inp_feat(196), I5 =>  inp_feat(373)); 
C_35_S_0_L_5_inst : LUT6 generic map(INIT => "0100011111111010001001111111101100001110111110110010000111011101") port map( O =>C_35_S_0_L_5_out, I0 =>  inp_feat(162), I1 =>  inp_feat(393), I2 =>  inp_feat(39), I3 =>  inp_feat(312), I4 =>  inp_feat(166), I5 =>  inp_feat(82)); 
C_35_S_1_L_0_inst : LUT6 generic map(INIT => "1111100110110010000000100000110000000000000000100011111000010000") port map( O =>C_35_S_1_L_0_out, I0 =>  inp_feat(493), I1 =>  inp_feat(429), I2 =>  inp_feat(226), I3 =>  inp_feat(162), I4 =>  inp_feat(280), I5 =>  inp_feat(321)); 
C_35_S_1_L_1_inst : LUT6 generic map(INIT => "1100011011111010111111101010001000000011101100001011000000000000") port map( O =>C_35_S_1_L_1_out, I0 =>  inp_feat(162), I1 =>  inp_feat(91), I2 =>  inp_feat(360), I3 =>  inp_feat(214), I4 =>  inp_feat(17), I5 =>  inp_feat(307)); 
C_35_S_1_L_2_inst : LUT6 generic map(INIT => "1011001110111000100001101111101001110110111000110000110111010100") port map( O =>C_35_S_1_L_2_out, I0 =>  inp_feat(162), I1 =>  inp_feat(235), I2 =>  inp_feat(394), I3 =>  inp_feat(264), I4 =>  inp_feat(468), I5 =>  inp_feat(4)); 
C_35_S_1_L_3_inst : LUT6 generic map(INIT => "1111100011111100011001000110010000000000000101001111010000110000") port map( O =>C_35_S_1_L_3_out, I0 =>  inp_feat(185), I1 =>  inp_feat(177), I2 =>  inp_feat(166), I3 =>  inp_feat(320), I4 =>  inp_feat(196), I5 =>  inp_feat(373)); 
C_35_S_1_L_4_inst : LUT6 generic map(INIT => "0100011111111010001001111111101100001110111110110010000111011101") port map( O =>C_35_S_1_L_4_out, I0 =>  inp_feat(162), I1 =>  inp_feat(393), I2 =>  inp_feat(39), I3 =>  inp_feat(312), I4 =>  inp_feat(166), I5 =>  inp_feat(82)); 
C_35_S_1_L_5_inst : LUT6 generic map(INIT => "1111011010110010000101010010111111100111000001110100110000101100") port map( O =>C_35_S_1_L_5_out, I0 =>  inp_feat(393), I1 =>  inp_feat(288), I2 =>  inp_feat(179), I3 =>  inp_feat(242), I4 =>  inp_feat(166), I5 =>  inp_feat(82)); 
C_35_S_2_L_0_inst : LUT6 generic map(INIT => "0111011111110110111111100010100000000110101000001000000000000000") port map( O =>C_35_S_2_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(278), I2 =>  inp_feat(166), I3 =>  inp_feat(214), I4 =>  inp_feat(17), I5 =>  inp_feat(307)); 
C_35_S_2_L_1_inst : LUT6 generic map(INIT => "1111100110111101111110000110110100000001100101110001000010000010") port map( O =>C_35_S_2_L_1_out, I0 =>  inp_feat(361), I1 =>  inp_feat(254), I2 =>  inp_feat(245), I3 =>  inp_feat(490), I4 =>  inp_feat(119), I5 =>  inp_feat(500)); 
C_35_S_2_L_2_inst : LUT6 generic map(INIT => "1110101011100100110011111111010100101110111011001111111111011010") port map( O =>C_35_S_2_L_2_out, I0 =>  inp_feat(61), I1 =>  inp_feat(13), I2 =>  inp_feat(343), I3 =>  inp_feat(178), I4 =>  inp_feat(478), I5 =>  inp_feat(476)); 
C_35_S_2_L_3_inst : LUT6 generic map(INIT => "1011001011011011101100100011111101010111010110010001010000000000") port map( O =>C_35_S_2_L_3_out, I0 =>  inp_feat(296), I1 =>  inp_feat(473), I2 =>  inp_feat(426), I3 =>  inp_feat(202), I4 =>  inp_feat(17), I5 =>  inp_feat(307)); 
C_35_S_2_L_4_inst : LUT6 generic map(INIT => "0001101111001001101011000001000000110010001110110011111000100010") port map( O =>C_35_S_2_L_4_out, I0 =>  inp_feat(307), I1 =>  inp_feat(292), I2 =>  inp_feat(507), I3 =>  inp_feat(245), I4 =>  inp_feat(360), I5 =>  inp_feat(130)); 
C_35_S_2_L_5_inst : LUT6 generic map(INIT => "0001111110001111101101110000111011001111010011110000000100001001") port map( O =>C_35_S_2_L_5_out, I0 =>  inp_feat(395), I1 =>  inp_feat(500), I2 =>  inp_feat(226), I3 =>  inp_feat(166), I4 =>  inp_feat(177), I5 =>  inp_feat(255)); 
C_35_S_3_L_0_inst : LUT6 generic map(INIT => "1100110011011010010000000011111110000000100100101000000010001010") port map( O =>C_35_S_3_L_0_out, I0 =>  inp_feat(321), I1 =>  inp_feat(81), I2 =>  inp_feat(468), I3 =>  inp_feat(230), I4 =>  inp_feat(177), I5 =>  inp_feat(255)); 
C_35_S_3_L_1_inst : LUT6 generic map(INIT => "0110011011111010111010000110001000100000111100001000000011110000") port map( O =>C_35_S_3_L_1_out, I0 =>  inp_feat(214), I1 =>  inp_feat(257), I2 =>  inp_feat(307), I3 =>  inp_feat(434), I4 =>  inp_feat(46), I5 =>  inp_feat(162)); 
C_35_S_3_L_2_inst : LUT6 generic map(INIT => "1111101111001011100011001001000000110010101110110011111000100010") port map( O =>C_35_S_3_L_2_out, I0 =>  inp_feat(307), I1 =>  inp_feat(292), I2 =>  inp_feat(507), I3 =>  inp_feat(245), I4 =>  inp_feat(360), I5 =>  inp_feat(130)); 
C_35_S_3_L_3_inst : LUT6 generic map(INIT => "0010111100010011100100100000001001010011100000101100000000000000") port map( O =>C_35_S_3_L_3_out, I0 =>  inp_feat(500), I1 =>  inp_feat(226), I2 =>  inp_feat(177), I3 =>  inp_feat(166), I4 =>  inp_feat(280), I5 =>  inp_feat(367)); 
C_35_S_3_L_4_inst : LUT6 generic map(INIT => "1101101100010011011110100000101010110010011000100010100010100000") port map( O =>C_35_S_3_L_4_out, I0 =>  inp_feat(465), I1 =>  inp_feat(429), I2 =>  inp_feat(488), I3 =>  inp_feat(229), I4 =>  inp_feat(330), I5 =>  inp_feat(124)); 
C_35_S_3_L_5_inst : LUT6 generic map(INIT => "1100001001110000000101100111100000000001000100011110111011100000") port map( O =>C_35_S_3_L_5_out, I0 =>  inp_feat(12), I1 =>  inp_feat(423), I2 =>  inp_feat(355), I3 =>  inp_feat(233), I4 =>  inp_feat(443), I5 =>  inp_feat(9)); 
C_35_S_4_L_0_inst : LUT6 generic map(INIT => "0000001010001111101001100000111001001111010011110000000000001001") port map( O =>C_35_S_4_L_0_out, I0 =>  inp_feat(395), I1 =>  inp_feat(500), I2 =>  inp_feat(226), I3 =>  inp_feat(166), I4 =>  inp_feat(177), I5 =>  inp_feat(255)); 
C_35_S_4_L_1_inst : LUT6 generic map(INIT => "1011100011110001110100001000000010010100100100100011001000110000") port map( O =>C_35_S_4_L_1_out, I0 =>  inp_feat(500), I1 =>  inp_feat(292), I2 =>  inp_feat(214), I3 =>  inp_feat(166), I4 =>  inp_feat(177), I5 =>  inp_feat(255)); 
C_35_S_4_L_2_inst : LUT6 generic map(INIT => "0110111001001010111010000110001000000000111100001000000011110000") port map( O =>C_35_S_4_L_2_out, I0 =>  inp_feat(214), I1 =>  inp_feat(257), I2 =>  inp_feat(307), I3 =>  inp_feat(434), I4 =>  inp_feat(46), I5 =>  inp_feat(162)); 
C_35_S_4_L_3_inst : LUT6 generic map(INIT => "1101001010010101101111101001110110010110111101000000000010000000") port map( O =>C_35_S_4_L_3_out, I0 =>  inp_feat(15), I1 =>  inp_feat(486), I2 =>  inp_feat(175), I3 =>  inp_feat(234), I4 =>  inp_feat(17), I5 =>  inp_feat(307)); 
C_35_S_4_L_4_inst : LUT6 generic map(INIT => "1101011010000100101011110000010000000111000000110000100100000000") port map( O =>C_35_S_4_L_4_out, I0 =>  inp_feat(360), I1 =>  inp_feat(278), I2 =>  inp_feat(413), I3 =>  inp_feat(166), I4 =>  inp_feat(468), I5 =>  inp_feat(151)); 
C_35_S_4_L_5_inst : LUT6 generic map(INIT => "0000111110001010110011100000110010000001010000010000101000000011") port map( O =>C_35_S_4_L_5_out, I0 =>  inp_feat(17), I1 =>  inp_feat(82), I2 =>  inp_feat(318), I3 =>  inp_feat(93), I4 =>  inp_feat(278), I5 =>  inp_feat(135)); 
C_35_S_5_L_0_inst : LUT6 generic map(INIT => "1001111101100100100111111100000000000000000000000010100000000000") port map( O =>C_35_S_5_L_0_out, I0 =>  inp_feat(500), I1 =>  inp_feat(17), I2 =>  inp_feat(278), I3 =>  inp_feat(307), I4 =>  inp_feat(224), I5 =>  inp_feat(378)); 
C_35_S_5_L_1_inst : LUT6 generic map(INIT => "0010001000000000111111111110110000100000001000001111111011000000") port map( O =>C_35_S_5_L_1_out, I0 =>  inp_feat(373), I1 =>  inp_feat(219), I2 =>  inp_feat(123), I3 =>  inp_feat(59), I4 =>  inp_feat(187), I5 =>  inp_feat(9)); 
C_35_S_5_L_2_inst : LUT6 generic map(INIT => "1110001001110000110111100111100000000001000100011110111011100000") port map( O =>C_35_S_5_L_2_out, I0 =>  inp_feat(12), I1 =>  inp_feat(423), I2 =>  inp_feat(355), I3 =>  inp_feat(233), I4 =>  inp_feat(443), I5 =>  inp_feat(9)); 
C_35_S_5_L_3_inst : LUT6 generic map(INIT => "0110110001011100010110101111110100000000010011001100100001110100") port map( O =>C_35_S_5_L_3_out, I0 =>  inp_feat(226), I1 =>  inp_feat(359), I2 =>  inp_feat(330), I3 =>  inp_feat(429), I4 =>  inp_feat(428), I5 =>  inp_feat(408)); 
C_35_S_5_L_4_inst : LUT6 generic map(INIT => "1011110110011101100111010000001110011101000100010011111100000001") port map( O =>C_35_S_5_L_4_out, I0 =>  inp_feat(321), I1 =>  inp_feat(180), I2 =>  inp_feat(344), I3 =>  inp_feat(11), I4 =>  inp_feat(422), I5 =>  inp_feat(283)); 
C_35_S_5_L_5_inst : LUT6 generic map(INIT => "0010010010100000110110001111110100000111000010000010101011111110") port map( O =>C_35_S_5_L_5_out, I0 =>  inp_feat(176), I1 =>  inp_feat(166), I2 =>  inp_feat(278), I3 =>  inp_feat(143), I4 =>  inp_feat(341), I5 =>  inp_feat(408)); 
C_36_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111010111111101111100011111100111110001000100010000000") port map( O =>C_36_S_0_L_0_out, I0 =>  inp_feat(195), I1 =>  inp_feat(48), I2 =>  inp_feat(426), I3 =>  inp_feat(385), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_36_S_0_L_1_inst : LUT6 generic map(INIT => "1111111111111101111110011010110011111101100100010100010001010100") port map( O =>C_36_S_0_L_1_out, I0 =>  inp_feat(186), I1 =>  inp_feat(458), I2 =>  inp_feat(482), I3 =>  inp_feat(440), I4 =>  inp_feat(456), I5 =>  inp_feat(232)); 
C_36_S_0_L_2_inst : LUT6 generic map(INIT => "1110111001001000111111111111111001101000110010001111111011100000") port map( O =>C_36_S_0_L_2_out, I0 =>  inp_feat(150), I1 =>  inp_feat(90), I2 =>  inp_feat(230), I3 =>  inp_feat(383), I4 =>  inp_feat(455), I5 =>  inp_feat(64)); 
C_36_S_0_L_3_inst : LUT6 generic map(INIT => "1110101101001010111111101111110011111000111000000110000000000000") port map( O =>C_36_S_0_L_3_out, I0 =>  inp_feat(90), I1 =>  inp_feat(48), I2 =>  inp_feat(426), I3 =>  inp_feat(64), I4 =>  inp_feat(262), I5 =>  inp_feat(9)); 
C_36_S_0_L_4_inst : LUT6 generic map(INIT => "1110111001101000111111011110101001111110001010001110101011101000") port map( O =>C_36_S_0_L_4_out, I0 =>  inp_feat(317), I1 =>  inp_feat(90), I2 =>  inp_feat(335), I3 =>  inp_feat(214), I4 =>  inp_feat(407), I5 =>  inp_feat(25)); 
C_36_S_0_L_5_inst : LUT6 generic map(INIT => "0110110101011110111011101110000011111111111010101111111011101001") port map( O =>C_36_S_0_L_5_out, I0 =>  inp_feat(82), I1 =>  inp_feat(465), I2 =>  inp_feat(80), I3 =>  inp_feat(457), I4 =>  inp_feat(168), I5 =>  inp_feat(290)); 
C_36_S_1_L_0_inst : LUT6 generic map(INIT => "1110111111001111111111111010100110001111000001111111101100000000") port map( O =>C_36_S_1_L_0_out, I0 =>  inp_feat(65), I1 =>  inp_feat(84), I2 =>  inp_feat(139), I3 =>  inp_feat(457), I4 =>  inp_feat(166), I5 =>  inp_feat(64)); 
C_36_S_1_L_1_inst : LUT6 generic map(INIT => "1111110011101000111111001000100001010110100011001111111010101000") port map( O =>C_36_S_1_L_1_out, I0 =>  inp_feat(224), I1 =>  inp_feat(383), I2 =>  inp_feat(385), I3 =>  inp_feat(150), I4 =>  inp_feat(120), I5 =>  inp_feat(199)); 
C_36_S_1_L_2_inst : LUT6 generic map(INIT => "1111000011101110111111101111110011101000111111100111000011101000") port map( O =>C_36_S_1_L_2_out, I0 =>  inp_feat(317), I1 =>  inp_feat(458), I2 =>  inp_feat(150), I3 =>  inp_feat(354), I4 =>  inp_feat(186), I5 =>  inp_feat(167)); 
C_36_S_1_L_3_inst : LUT6 generic map(INIT => "1110110010000000111011101010100011101000100000000000100010100000") port map( O =>C_36_S_1_L_3_out, I0 =>  inp_feat(426), I1 =>  inp_feat(177), I2 =>  inp_feat(473), I3 =>  inp_feat(16), I4 =>  inp_feat(218), I5 =>  inp_feat(196)); 
C_36_S_1_L_4_inst : LUT6 generic map(INIT => "0110100011100100111000001111111011111110111111111110110011111101") port map( O =>C_36_S_1_L_4_out, I0 =>  inp_feat(317), I1 =>  inp_feat(232), I2 =>  inp_feat(440), I3 =>  inp_feat(413), I4 =>  inp_feat(476), I5 =>  inp_feat(168)); 
C_36_S_1_L_5_inst : LUT6 generic map(INIT => "1000111011100110010011101111100011101111101010001110111010100000") port map( O =>C_36_S_1_L_5_out, I0 =>  inp_feat(482), I1 =>  inp_feat(232), I2 =>  inp_feat(164), I3 =>  inp_feat(343), I4 =>  inp_feat(346), I5 =>  inp_feat(319)); 
C_36_S_2_L_0_inst : LUT6 generic map(INIT => "1110111111101110111111111110001010010000110010001111111010001000") port map( O =>C_36_S_2_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(458), I2 =>  inp_feat(237), I3 =>  inp_feat(50), I4 =>  inp_feat(319), I5 =>  inp_feat(150)); 
C_36_S_2_L_1_inst : LUT6 generic map(INIT => "1110111011101000111111111111101001111100111010001111111111111110") port map( O =>C_36_S_2_L_1_out, I0 =>  inp_feat(473), I1 =>  inp_feat(458), I2 =>  inp_feat(264), I3 =>  inp_feat(48), I4 =>  inp_feat(407), I5 =>  inp_feat(303)); 
C_36_S_2_L_2_inst : LUT6 generic map(INIT => "1110001011101010111111111010101000110011101010101011111110101010") port map( O =>C_36_S_2_L_2_out, I0 =>  inp_feat(426), I1 =>  inp_feat(170), I2 =>  inp_feat(451), I3 =>  inp_feat(446), I4 =>  inp_feat(74), I5 =>  inp_feat(32)); 
C_36_S_2_L_3_inst : LUT6 generic map(INIT => "1111110111100000010111101110111011101100100010001110111011101100") port map( O =>C_36_S_2_L_3_out, I0 =>  inp_feat(315), I1 =>  inp_feat(426), I2 =>  inp_feat(48), I3 =>  inp_feat(232), I4 =>  inp_feat(489), I5 =>  inp_feat(446)); 
C_36_S_2_L_4_inst : LUT6 generic map(INIT => "0110010111111110111111111111111111111111111111001111111111111110") port map( O =>C_36_S_2_L_4_out, I0 =>  inp_feat(126), I1 =>  inp_feat(167), I2 =>  inp_feat(237), I3 =>  inp_feat(168), I4 =>  inp_feat(290), I5 =>  inp_feat(139)); 
C_36_S_2_L_5_inst : LUT6 generic map(INIT => "1111110111010000111011111111111011111111111111011111111111111000") port map( O =>C_36_S_2_L_5_out, I0 =>  inp_feat(471), I1 =>  inp_feat(426), I2 =>  inp_feat(482), I3 =>  inp_feat(176), I4 =>  inp_feat(170), I5 =>  inp_feat(453)); 
C_36_S_3_L_0_inst : LUT6 generic map(INIT => "1111111110101111111111110010111111111111100011000111111100101100") port map( O =>C_36_S_3_L_0_out, I0 =>  inp_feat(482), I1 =>  inp_feat(222), I2 =>  inp_feat(74), I3 =>  inp_feat(150), I4 =>  inp_feat(456), I5 =>  inp_feat(32)); 
C_36_S_3_L_1_inst : LUT6 generic map(INIT => "0011001011111110111110101011101011111011111110101111101010111010") port map( O =>C_36_S_3_L_1_out, I0 =>  inp_feat(482), I1 =>  inp_feat(435), I2 =>  inp_feat(458), I3 =>  inp_feat(354), I4 =>  inp_feat(446), I5 =>  inp_feat(453)); 
C_36_S_3_L_2_inst : LUT6 generic map(INIT => "1110111101100010111111101111000011110010001000001011001001000000") port map( O =>C_36_S_3_L_2_out, I0 =>  inp_feat(497), I1 =>  inp_feat(24), I2 =>  inp_feat(237), I3 =>  inp_feat(383), I4 =>  inp_feat(422), I5 =>  inp_feat(167)); 
C_36_S_3_L_3_inst : LUT6 generic map(INIT => "1111001010101000111111111110010011011100000000001010000011000000") port map( O =>C_36_S_3_L_3_out, I0 =>  inp_feat(482), I1 =>  inp_feat(383), I2 =>  inp_feat(344), I3 =>  inp_feat(426), I4 =>  inp_feat(369), I5 =>  inp_feat(457)); 
C_36_S_3_L_4_inst : LUT6 generic map(INIT => "1101111111110111000111111111110111111111111111111111111111011100") port map( O =>C_36_S_3_L_4_out, I0 =>  inp_feat(389), I1 =>  inp_feat(264), I2 =>  inp_feat(89), I3 =>  inp_feat(95), I4 =>  inp_feat(456), I5 =>  inp_feat(290)); 
C_36_S_3_L_5_inst : LUT6 generic map(INIT => "1000111010111111111111111111011111111111111011000011111111001100") port map( O =>C_36_S_3_L_5_out, I0 =>  inp_feat(458), I1 =>  inp_feat(171), I2 =>  inp_feat(300), I3 =>  inp_feat(493), I4 =>  inp_feat(130), I5 =>  inp_feat(461)); 
C_36_S_4_L_0_inst : LUT6 generic map(INIT => "1110100011111110111111000110101001001000100000101100000010000000") port map( O =>C_36_S_4_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(90), I2 =>  inp_feat(224), I3 =>  inp_feat(244), I4 =>  inp_feat(167), I5 =>  inp_feat(271)); 
C_36_S_4_L_1_inst : LUT6 generic map(INIT => "1011110001010100111111011111000110010100110100001101010011010000") port map( O =>C_36_S_4_L_1_out, I0 =>  inp_feat(449), I1 =>  inp_feat(237), I2 =>  inp_feat(66), I3 =>  inp_feat(7), I4 =>  inp_feat(332), I5 =>  inp_feat(64)); 
C_36_S_4_L_2_inst : LUT6 generic map(INIT => "1110110011111110111111111111000000101000101000001111111010101000") port map( O =>C_36_S_4_L_2_out, I0 =>  inp_feat(264), I1 =>  inp_feat(237), I2 =>  inp_feat(368), I3 =>  inp_feat(24), I4 =>  inp_feat(325), I5 =>  inp_feat(64)); 
C_36_S_4_L_3_inst : LUT6 generic map(INIT => "1110111011100111111111111101111111111111111111110100111101111110") port map( O =>C_36_S_4_L_3_out, I0 =>  inp_feat(317), I1 =>  inp_feat(167), I2 =>  inp_feat(111), I3 =>  inp_feat(72), I4 =>  inp_feat(130), I5 =>  inp_feat(461)); 
C_36_S_4_L_4_inst : LUT6 generic map(INIT => "0001101000101000100110110010101011111110101010101011101000001000") port map( O =>C_36_S_4_L_4_out, I0 =>  inp_feat(426), I1 =>  inp_feat(306), I2 =>  inp_feat(321), I3 =>  inp_feat(177), I4 =>  inp_feat(333), I5 =>  inp_feat(493)); 
C_36_S_4_L_5_inst : LUT6 generic map(INIT => "1011110011100110111111111111011101110000111011001111110111111111") port map( O =>C_36_S_4_L_5_out, I0 =>  inp_feat(243), I1 =>  inp_feat(171), I2 =>  inp_feat(426), I3 =>  inp_feat(174), I4 =>  inp_feat(170), I5 =>  inp_feat(156)); 
C_36_S_5_L_0_inst : LUT6 generic map(INIT => "0010111100001111111111111111111011101111000011111101011111111111") port map( O =>C_36_S_5_L_0_out, I0 =>  inp_feat(448), I1 =>  inp_feat(0), I2 =>  inp_feat(160), I3 =>  inp_feat(383), I4 =>  inp_feat(399), I5 =>  inp_feat(381)); 
C_36_S_5_L_1_inst : LUT6 generic map(INIT => "1110100011001110111111101110100001101000111010001110111011101000") port map( O =>C_36_S_5_L_1_out, I0 =>  inp_feat(482), I1 =>  inp_feat(237), I2 =>  inp_feat(335), I3 =>  inp_feat(79), I4 =>  inp_feat(407), I5 =>  inp_feat(381)); 
C_36_S_5_L_2_inst : LUT6 generic map(INIT => "1111111111111000101011001010100001101110101101001111101010000000") port map( O =>C_36_S_5_L_2_out, I0 =>  inp_feat(426), I1 =>  inp_feat(232), I2 =>  inp_feat(195), I3 =>  inp_feat(335), I4 =>  inp_feat(81), I5 =>  inp_feat(489)); 
C_36_S_5_L_3_inst : LUT6 generic map(INIT => "0100101011001110111111101111111111100100111011001110111000101110") port map( O =>C_36_S_5_L_3_out, I0 =>  inp_feat(482), I1 =>  inp_feat(458), I2 =>  inp_feat(317), I3 =>  inp_feat(470), I4 =>  inp_feat(157), I5 =>  inp_feat(37)); 
C_36_S_5_L_4_inst : LUT6 generic map(INIT => "1111111111100111111111101111111111111111111100011101011111110011") port map( O =>C_36_S_5_L_4_out, I0 =>  inp_feat(59), I1 =>  inp_feat(11), I2 =>  inp_feat(90), I3 =>  inp_feat(346), I4 =>  inp_feat(29), I5 =>  inp_feat(457)); 
C_36_S_5_L_5_inst : LUT6 generic map(INIT => "1100111011111111100000001110100011111011010111111111111010101100") port map( O =>C_36_S_5_L_5_out, I0 =>  inp_feat(84), I1 =>  inp_feat(383), I2 =>  inp_feat(66), I3 =>  inp_feat(93), I4 =>  inp_feat(458), I5 =>  inp_feat(343)); 
C_37_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000010000011100000011000001110011011101111111") port map( O =>C_37_S_0_L_0_out, I0 =>  inp_feat(195), I1 =>  inp_feat(48), I2 =>  inp_feat(426), I3 =>  inp_feat(385), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_0_L_1_inst : LUT6 generic map(INIT => "1100000100000111000100110001111110100011000001111111111101011111") port map( O =>C_37_S_0_L_1_out, I0 =>  inp_feat(150), I1 =>  inp_feat(230), I2 =>  inp_feat(232), I3 =>  inp_feat(386), I4 =>  inp_feat(383), I5 =>  inp_feat(246)); 
C_37_S_0_L_2_inst : LUT6 generic map(INIT => "1111101011110011010101001111111111000000110000100000010000000000") port map( O =>C_37_S_0_L_2_out, I0 =>  inp_feat(7), I1 =>  inp_feat(245), I2 =>  inp_feat(199), I3 =>  inp_feat(383), I4 =>  inp_feat(372), I5 =>  inp_feat(266)); 
C_37_S_0_L_3_inst : LUT6 generic map(INIT => "0000100000000010000000001001101011001010000110100010101101111111") port map( O =>C_37_S_0_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(335), I2 =>  inp_feat(90), I3 =>  inp_feat(66), I4 =>  inp_feat(385), I5 =>  inp_feat(383)); 
C_37_S_0_L_4_inst : LUT6 generic map(INIT => "1010111100010111001100110101011100000000000000110000000000000000") port map( O =>C_37_S_0_L_4_out, I0 =>  inp_feat(150), I1 =>  inp_feat(232), I2 =>  inp_feat(458), I3 =>  inp_feat(315), I4 =>  inp_feat(372), I5 =>  inp_feat(432)); 
C_37_S_0_L_5_inst : LUT6 generic map(INIT => "0010011100100101110011000000010100000101010001110011011101111111") port map( O =>C_37_S_0_L_5_out, I0 =>  inp_feat(482), I1 =>  inp_feat(385), I2 =>  inp_feat(458), I3 =>  inp_feat(237), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_37_S_1_L_0_inst : LUT6 generic map(INIT => "1100000100000111000100110001111110100011000001111111111101011111") port map( O =>C_37_S_1_L_0_out, I0 =>  inp_feat(150), I1 =>  inp_feat(230), I2 =>  inp_feat(232), I3 =>  inp_feat(386), I4 =>  inp_feat(383), I5 =>  inp_feat(246)); 
C_37_S_1_L_1_inst : LUT6 generic map(INIT => "1111101011110011010101001111111111000000110000100000010000000000") port map( O =>C_37_S_1_L_1_out, I0 =>  inp_feat(7), I1 =>  inp_feat(245), I2 =>  inp_feat(199), I3 =>  inp_feat(383), I4 =>  inp_feat(372), I5 =>  inp_feat(266)); 
C_37_S_1_L_2_inst : LUT6 generic map(INIT => "0000100000000010000000001001101011001010000110100010101101111111") port map( O =>C_37_S_1_L_2_out, I0 =>  inp_feat(100), I1 =>  inp_feat(335), I2 =>  inp_feat(90), I3 =>  inp_feat(66), I4 =>  inp_feat(385), I5 =>  inp_feat(383)); 
C_37_S_1_L_3_inst : LUT6 generic map(INIT => "1010111100010111001100110101011100000000000000110000000000000000") port map( O =>C_37_S_1_L_3_out, I0 =>  inp_feat(150), I1 =>  inp_feat(232), I2 =>  inp_feat(458), I3 =>  inp_feat(315), I4 =>  inp_feat(372), I5 =>  inp_feat(432)); 
C_37_S_1_L_4_inst : LUT6 generic map(INIT => "0010011100100101110011000000010100000101010001110011011101111111") port map( O =>C_37_S_1_L_4_out, I0 =>  inp_feat(482), I1 =>  inp_feat(385), I2 =>  inp_feat(458), I3 =>  inp_feat(237), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_37_S_1_L_5_inst : LUT6 generic map(INIT => "1000101010100000010001000000000011010110111010001111010001110100") port map( O =>C_37_S_1_L_5_out, I0 =>  inp_feat(463), I1 =>  inp_feat(488), I2 =>  inp_feat(104), I3 =>  inp_feat(312), I4 =>  inp_feat(482), I5 =>  inp_feat(232)); 
C_37_S_2_L_0_inst : LUT6 generic map(INIT => "0000101010000000001011000000000011100110111110001111110011110100") port map( O =>C_37_S_2_L_0_out, I0 =>  inp_feat(224), I1 =>  inp_feat(488), I2 =>  inp_feat(104), I3 =>  inp_feat(312), I4 =>  inp_feat(482), I5 =>  inp_feat(232)); 
C_37_S_2_L_1_inst : LUT6 generic map(INIT => "1110001100010011000100110111011100000111000001010000000100000111") port map( O =>C_37_S_2_L_1_out, I0 =>  inp_feat(317), I1 =>  inp_feat(232), I2 =>  inp_feat(482), I3 =>  inp_feat(335), I4 =>  inp_feat(372), I5 =>  inp_feat(221)); 
C_37_S_2_L_2_inst : LUT6 generic map(INIT => "1101010110001100111111110000011010001000000001001000000000001100") port map( O =>C_37_S_2_L_2_out, I0 =>  inp_feat(427), I1 =>  inp_feat(301), I2 =>  inp_feat(415), I3 =>  inp_feat(287), I4 =>  inp_feat(484), I5 =>  inp_feat(42)); 
C_37_S_2_L_3_inst : LUT6 generic map(INIT => "0000000001000001000000010011011100000001010100110001111101111111") port map( O =>C_37_S_2_L_3_out, I0 =>  inp_feat(317), I1 =>  inp_feat(458), I2 =>  inp_feat(456), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_2_L_4_inst : LUT6 generic map(INIT => "1001101001010111110011001101100000000000101011100001000110000000") port map( O =>C_37_S_2_L_4_out, I0 =>  inp_feat(456), I1 =>  inp_feat(317), I2 =>  inp_feat(441), I3 =>  inp_feat(28), I4 =>  inp_feat(436), I5 =>  inp_feat(104)); 
C_37_S_2_L_5_inst : LUT6 generic map(INIT => "1011000100010111100101010111111100000001000110111001011101011111") port map( O =>C_37_S_2_L_5_out, I0 =>  inp_feat(463), I1 =>  inp_feat(458), I2 =>  inp_feat(426), I3 =>  inp_feat(315), I4 =>  inp_feat(380), I5 =>  inp_feat(202)); 
C_37_S_3_L_0_inst : LUT6 generic map(INIT => "0000000100010001100110110000000000010011000000000111111100000001") port map( O =>C_37_S_3_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(458), I2 =>  inp_feat(246), I3 =>  inp_feat(204), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_3_L_1_inst : LUT6 generic map(INIT => "1000001111000111000001110010001001100000000000000000000000000000") port map( O =>C_37_S_3_L_1_out, I0 =>  inp_feat(441), I1 =>  inp_feat(183), I2 =>  inp_feat(413), I3 =>  inp_feat(482), I4 =>  inp_feat(74), I5 =>  inp_feat(366)); 
C_37_S_3_L_2_inst : LUT6 generic map(INIT => "1100111111011010110011101100111000000111000000110000110010011001") port map( O =>C_37_S_3_L_2_out, I0 =>  inp_feat(26), I1 =>  inp_feat(35), I2 =>  inp_feat(215), I3 =>  inp_feat(365), I4 =>  inp_feat(353), I5 =>  inp_feat(42)); 
C_37_S_3_L_3_inst : LUT6 generic map(INIT => "1100010001010101000011010111111100000001000101010001011101011111") port map( O =>C_37_S_3_L_3_out, I0 =>  inp_feat(232), I1 =>  inp_feat(176), I2 =>  inp_feat(66), I3 =>  inp_feat(317), I4 =>  inp_feat(383), I5 =>  inp_feat(202)); 
C_37_S_3_L_4_inst : LUT6 generic map(INIT => "0001010111101111110111101110100000000110111110000110000010000000") port map( O =>C_37_S_3_L_4_out, I0 =>  inp_feat(226), I1 =>  inp_feat(489), I2 =>  inp_feat(334), I3 =>  inp_feat(7), I4 =>  inp_feat(431), I5 =>  inp_feat(161)); 
C_37_S_3_L_5_inst : LUT6 generic map(INIT => "1000010100011111111011111100011100000000100000100001000000000000") port map( O =>C_37_S_3_L_5_out, I0 =>  inp_feat(322), I1 =>  inp_feat(45), I2 =>  inp_feat(458), I3 =>  inp_feat(482), I4 =>  inp_feat(289), I5 =>  inp_feat(266)); 
C_37_S_4_L_0_inst : LUT6 generic map(INIT => "0101000100110101010101110000000000110011001000000111111100000011") port map( O =>C_37_S_4_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(458), I2 =>  inp_feat(246), I3 =>  inp_feat(204), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_4_L_1_inst : LUT6 generic map(INIT => "1000101001010010100101001100110001111010001010000100110011001100") port map( O =>C_37_S_4_L_1_out, I0 =>  inp_feat(176), I1 =>  inp_feat(325), I2 =>  inp_feat(48), I3 =>  inp_feat(482), I4 =>  inp_feat(232), I5 =>  inp_feat(213)); 
C_37_S_4_L_2_inst : LUT6 generic map(INIT => "0000001110111000100110000010000011000100100101001010100010000000") port map( O =>C_37_S_4_L_2_out, I0 =>  inp_feat(203), I1 =>  inp_feat(211), I2 =>  inp_feat(470), I3 =>  inp_feat(403), I4 =>  inp_feat(177), I5 =>  inp_feat(315)); 
C_37_S_4_L_3_inst : LUT6 generic map(INIT => "1101000011000001101110010001111110001101111101110001011101111111") port map( O =>C_37_S_4_L_3_out, I0 =>  inp_feat(232), I1 =>  inp_feat(237), I2 =>  inp_feat(456), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_4_L_4_inst : LUT6 generic map(INIT => "0011100000001001000110110011011100101001110100010001111101111111") port map( O =>C_37_S_4_L_4_out, I0 =>  inp_feat(317), I1 =>  inp_feat(458), I2 =>  inp_feat(456), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_4_L_5_inst : LUT6 generic map(INIT => "1110010111100011000010101000010111101000000000100000110000000001") port map( O =>C_37_S_4_L_5_out, I0 =>  inp_feat(110), I1 =>  inp_feat(307), I2 =>  inp_feat(411), I3 =>  inp_feat(303), I4 =>  inp_feat(42), I5 =>  inp_feat(484)); 
C_37_S_5_L_0_inst : LUT6 generic map(INIT => "0001001000001000000110000100100000001000100011000000100010001110") port map( O =>C_37_S_5_L_0_out, I0 =>  inp_feat(108), I1 =>  inp_feat(102), I2 =>  inp_feat(90), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_5_L_1_inst : LUT6 generic map(INIT => "1101000000011101101000110001011110011011111111110001011101110111") port map( O =>C_37_S_5_L_1_out, I0 =>  inp_feat(150), I1 =>  inp_feat(90), I2 =>  inp_feat(468), I3 =>  inp_feat(482), I4 =>  inp_feat(213), I5 =>  inp_feat(232)); 
C_37_S_5_L_2_inst : LUT6 generic map(INIT => "1110111101011011111110110011001011111011001100000010000000000000") port map( O =>C_37_S_5_L_2_out, I0 =>  inp_feat(282), I1 =>  inp_feat(391), I2 =>  inp_feat(187), I3 =>  inp_feat(1), I4 =>  inp_feat(431), I5 =>  inp_feat(161)); 
C_37_S_5_L_3_inst : LUT6 generic map(INIT => "0011000001000001000110010011011100001001000100010001111101111111") port map( O =>C_37_S_5_L_3_out, I0 =>  inp_feat(317), I1 =>  inp_feat(458), I2 =>  inp_feat(456), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_37_S_5_L_4_inst : LUT6 generic map(INIT => "0110000000101000111010000000100011111000101010001110000000000000") port map( O =>C_37_S_5_L_4_out, I0 =>  inp_feat(289), I1 =>  inp_feat(482), I2 =>  inp_feat(502), I3 =>  inp_feat(391), I4 =>  inp_feat(76), I5 =>  inp_feat(141)); 
C_37_S_5_L_5_inst : LUT6 generic map(INIT => "1111111110000111000110111101011100000000100101010001010100010111") port map( O =>C_37_S_5_L_5_out, I0 =>  inp_feat(232), I1 =>  inp_feat(335), I2 =>  inp_feat(315), I3 =>  inp_feat(81), I4 =>  inp_feat(385), I5 =>  inp_feat(305)); 
C_38_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000000000000010001011100000000000101110001011101111111") port map( O =>C_38_S_0_L_0_out, I0 =>  inp_feat(385), I1 =>  inp_feat(317), I2 =>  inp_feat(48), I3 =>  inp_feat(237), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_38_S_0_L_1_inst : LUT6 generic map(INIT => "0101011110111011000000110010101111110110101011110000101100101011") port map( O =>C_38_S_0_L_1_out, I0 =>  inp_feat(455), I1 =>  inp_feat(458), I2 =>  inp_feat(426), I3 =>  inp_feat(150), I4 =>  inp_feat(212), I5 =>  inp_feat(7)); 
C_38_S_0_L_2_inst : LUT6 generic map(INIT => "0000001000101000111011111111001011111101111010001111111011110010") port map( O =>C_38_S_0_L_2_out, I0 =>  inp_feat(91), I1 =>  inp_feat(232), I2 =>  inp_feat(204), I3 =>  inp_feat(315), I4 =>  inp_feat(383), I5 =>  inp_feat(497)); 
C_38_S_0_L_3_inst : LUT6 generic map(INIT => "1110101110101110111111010010000100000000000000001100000100000100") port map( O =>C_38_S_0_L_3_out, I0 =>  inp_feat(385), I1 =>  inp_feat(123), I2 =>  inp_feat(459), I3 =>  inp_feat(151), I4 =>  inp_feat(214), I5 =>  inp_feat(147)); 
C_38_S_0_L_4_inst : LUT6 generic map(INIT => "0000000000111111001001010101111100100010011111110011011101111111") port map( O =>C_38_S_0_L_4_out, I0 =>  inp_feat(237), I1 =>  inp_feat(468), I2 =>  inp_feat(482), I3 =>  inp_feat(458), I4 =>  inp_feat(66), I5 =>  inp_feat(473)); 
C_38_S_0_L_5_inst : LUT6 generic map(INIT => "1111111111100011111111111100001100001101010001000000010000000000") port map( O =>C_38_S_0_L_5_out, I0 =>  inp_feat(473), I1 =>  inp_feat(383), I2 =>  inp_feat(66), I3 =>  inp_feat(93), I4 =>  inp_feat(87), I5 =>  inp_feat(51)); 
C_38_S_1_L_0_inst : LUT6 generic map(INIT => "1011001110111111000100110011011111101001111111110001101100111111") port map( O =>C_38_S_1_L_0_out, I0 =>  inp_feat(482), I1 =>  inp_feat(458), I2 =>  inp_feat(426), I3 =>  inp_feat(150), I4 =>  inp_feat(212), I5 =>  inp_feat(7)); 
C_38_S_1_L_1_inst : LUT6 generic map(INIT => "0011001100001001100101011100110101110111001111110010110111011111") port map( O =>C_38_S_1_L_1_out, I0 =>  inp_feat(373), I1 =>  inp_feat(497), I2 =>  inp_feat(482), I3 =>  inp_feat(177), I4 =>  inp_feat(426), I5 =>  inp_feat(7)); 
C_38_S_1_L_2_inst : LUT6 generic map(INIT => "0001000100010101100001011110000010010001100111010000001100000001") port map( O =>C_38_S_1_L_2_out, I0 =>  inp_feat(444), I1 =>  inp_feat(28), I2 =>  inp_feat(359), I3 =>  inp_feat(383), I4 =>  inp_feat(150), I5 =>  inp_feat(194)); 
C_38_S_1_L_3_inst : LUT6 generic map(INIT => "0000110111000111000000011101111100001011100101110001011100111111") port map( O =>C_38_S_1_L_3_out, I0 =>  inp_feat(440), I1 =>  inp_feat(48), I2 =>  inp_feat(458), I3 =>  inp_feat(482), I4 =>  inp_feat(426), I5 =>  inp_feat(463)); 
C_38_S_1_L_4_inst : LUT6 generic map(INIT => "1001010111111101110101010011111111011101110111111101110101111111") port map( O =>C_38_S_1_L_4_out, I0 =>  inp_feat(90), I1 =>  inp_feat(385), I2 =>  inp_feat(66), I3 =>  inp_feat(386), I4 =>  inp_feat(383), I5 =>  inp_feat(2)); 
C_38_S_1_L_5_inst : LUT6 generic map(INIT => "1101001000001100111111101000110000001000001000101110111000001000") port map( O =>C_38_S_1_L_5_out, I0 =>  inp_feat(455), I1 =>  inp_feat(472), I2 =>  inp_feat(317), I3 =>  inp_feat(17), I4 =>  inp_feat(132), I5 =>  inp_feat(182)); 
C_38_S_2_L_0_inst : LUT6 generic map(INIT => "0010000100010101000100010101111111110001001110111111011101111111") port map( O =>C_38_S_2_L_0_out, I0 =>  inp_feat(317), I1 =>  inp_feat(232), I2 =>  inp_feat(48), I3 =>  inp_feat(150), I4 =>  inp_feat(383), I5 =>  inp_feat(456)); 
C_38_S_2_L_1_inst : LUT6 generic map(INIT => "1010001100000000010111110100110100111011000010010111111110001111") port map( O =>C_38_S_2_L_1_out, I0 =>  inp_feat(150), I1 =>  inp_feat(84), I2 =>  inp_feat(468), I3 =>  inp_feat(183), I4 =>  inp_feat(66), I5 =>  inp_feat(473)); 
C_38_S_2_L_2_inst : LUT6 generic map(INIT => "0011011100001101111000011011011111000111100101111101011101111111") port map( O =>C_38_S_2_L_2_out, I0 =>  inp_feat(90), I1 =>  inp_feat(458), I2 =>  inp_feat(317), I3 =>  inp_feat(232), I4 =>  inp_feat(66), I5 =>  inp_feat(473)); 
C_38_S_2_L_3_inst : LUT6 generic map(INIT => "1101000110011111110100111001100100010000000000000000000001000000") port map( O =>C_38_S_2_L_3_out, I0 =>  inp_feat(482), I1 =>  inp_feat(335), I2 =>  inp_feat(447), I3 =>  inp_feat(18), I4 =>  inp_feat(87), I5 =>  inp_feat(147)); 
C_38_S_2_L_4_inst : LUT6 generic map(INIT => "0000000000110000000100001111000000010001101100000111000011110010") port map( O =>C_38_S_2_L_4_out, I0 =>  inp_feat(245), I1 =>  inp_feat(456), I2 =>  inp_feat(51), I3 =>  inp_feat(232), I4 =>  inp_feat(150), I5 =>  inp_feat(64)); 
C_38_S_2_L_5_inst : LUT6 generic map(INIT => "0001100000000100000001010011111111111101010000010000000100000111") port map( O =>C_38_S_2_L_5_out, I0 =>  inp_feat(256), I1 =>  inp_feat(166), I2 =>  inp_feat(31), I3 =>  inp_feat(124), I4 =>  inp_feat(454), I5 =>  inp_feat(157)); 
C_38_S_3_L_0_inst : LUT6 generic map(INIT => "0010010100000111001100111001011111010001011101111111011111111111") port map( O =>C_38_S_3_L_0_out, I0 =>  inp_feat(195), I1 =>  inp_feat(426), I2 =>  inp_feat(385), I3 =>  inp_feat(232), I4 =>  inp_feat(66), I5 =>  inp_feat(473)); 
C_38_S_3_L_1_inst : LUT6 generic map(INIT => "1000000100011111001100000111101110011000011100001111101001110000") port map( O =>C_38_S_3_L_1_out, I0 =>  inp_feat(232), I1 =>  inp_feat(150), I2 =>  inp_feat(116), I3 =>  inp_feat(176), I4 =>  inp_feat(66), I5 =>  inp_feat(468)); 
C_38_S_3_L_2_inst : LUT6 generic map(INIT => "0101001100001001011100110111000101111101010100110100011111111111") port map( O =>C_38_S_3_L_2_out, I0 =>  inp_feat(317), I1 =>  inp_feat(232), I2 =>  inp_feat(385), I3 =>  inp_feat(48), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_38_S_3_L_3_inst : LUT6 generic map(INIT => "1101011000100010111100110010011011011010101000100001101010101010") port map( O =>C_38_S_3_L_3_out, I0 =>  inp_feat(160), I1 =>  inp_feat(232), I2 =>  inp_feat(385), I3 =>  inp_feat(48), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_38_S_3_L_4_inst : LUT6 generic map(INIT => "0000011100110101100101010011011101100101101101111111111101111111") port map( O =>C_38_S_3_L_4_out, I0 =>  inp_feat(458), I1 =>  inp_feat(150), I2 =>  inp_feat(385), I3 =>  inp_feat(176), I4 =>  inp_feat(468), I5 =>  inp_feat(66)); 
C_38_S_3_L_5_inst : LUT6 generic map(INIT => "1111110101000100111100001110100001110011111101111101000011110100") port map( O =>C_38_S_3_L_5_out, I0 =>  inp_feat(258), I1 =>  inp_feat(165), I2 =>  inp_feat(289), I3 =>  inp_feat(426), I4 =>  inp_feat(177), I5 =>  inp_feat(2)); 
C_38_S_4_L_0_inst : LUT6 generic map(INIT => "1111111000111011111111110001100111110111000000001111011100000000") port map( O =>C_38_S_4_L_0_out, I0 =>  inp_feat(335), I1 =>  inp_feat(214), I2 =>  inp_feat(173), I3 =>  inp_feat(325), I4 =>  inp_feat(150), I5 =>  inp_feat(64)); 
C_38_S_4_L_1_inst : LUT6 generic map(INIT => "0001101001011011010101110101101110011010001111010010111101110111") port map( O =>C_38_S_4_L_1_out, I0 =>  inp_feat(48), I1 =>  inp_feat(426), I2 =>  inp_feat(468), I3 =>  inp_feat(90), I4 =>  inp_feat(150), I5 =>  inp_feat(64)); 
C_38_S_4_L_2_inst : LUT6 generic map(INIT => "0001100100011101000110111111111111110011000100011111001100011001") port map( O =>C_38_S_4_L_2_out, I0 =>  inp_feat(458), I1 =>  inp_feat(482), I2 =>  inp_feat(2), I3 =>  inp_feat(106), I4 =>  inp_feat(226), I5 =>  inp_feat(199)); 
C_38_S_4_L_3_inst : LUT6 generic map(INIT => "1110100010001100111111101101001100010100000001001011010100000101") port map( O =>C_38_S_4_L_3_out, I0 =>  inp_feat(33), I1 =>  inp_feat(441), I2 =>  inp_feat(93), I3 =>  inp_feat(19), I4 =>  inp_feat(132), I5 =>  inp_feat(180)); 
C_38_S_4_L_4_inst : LUT6 generic map(INIT => "0001010101110100101100001111010111110000110100101011100111110001") port map( O =>C_38_S_4_L_4_out, I0 =>  inp_feat(383), I1 =>  inp_feat(456), I2 =>  inp_feat(378), I3 =>  inp_feat(463), I4 =>  inp_feat(66), I5 =>  inp_feat(258)); 
C_38_S_4_L_5_inst : LUT6 generic map(INIT => "1011101101011101100011010111011111101000001111110000110111111111") port map( O =>C_38_S_4_L_5_out, I0 =>  inp_feat(385), I1 =>  inp_feat(177), I2 =>  inp_feat(195), I3 =>  inp_feat(150), I4 =>  inp_feat(361), I5 =>  inp_feat(490)); 
C_38_S_5_L_0_inst : LUT6 generic map(INIT => "0001000100000001000100110101000110111001010101110100011111111111") port map( O =>C_38_S_5_L_0_out, I0 =>  inp_feat(317), I1 =>  inp_feat(232), I2 =>  inp_feat(385), I3 =>  inp_feat(48), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_38_S_5_L_1_inst : LUT6 generic map(INIT => "1001101110001101010110010101111101000111001100111001101101111111") port map( O =>C_38_S_5_L_1_out, I0 =>  inp_feat(317), I1 =>  inp_feat(90), I2 =>  inp_feat(456), I3 =>  inp_feat(383), I4 =>  inp_feat(150), I5 =>  inp_feat(64)); 
C_38_S_5_L_2_inst : LUT6 generic map(INIT => "0010001001011001000000110101111110000111001100111001101101111111") port map( O =>C_38_S_5_L_2_out, I0 =>  inp_feat(246), I1 =>  inp_feat(90), I2 =>  inp_feat(456), I3 =>  inp_feat(383), I4 =>  inp_feat(150), I5 =>  inp_feat(64)); 
C_38_S_5_L_3_inst : LUT6 generic map(INIT => "1001011011010101110011110000110000001100010011001111111111001100") port map( O =>C_38_S_5_L_3_out, I0 =>  inp_feat(216), I1 =>  inp_feat(61), I2 =>  inp_feat(426), I3 =>  inp_feat(383), I4 =>  inp_feat(473), I5 =>  inp_feat(66)); 
C_38_S_5_L_4_inst : LUT6 generic map(INIT => "0000100111100011101101010101111111100111100101111111011111111111") port map( O =>C_38_S_5_L_4_out, I0 =>  inp_feat(90), I1 =>  inp_feat(426), I2 =>  inp_feat(385), I3 =>  inp_feat(383), I4 =>  inp_feat(386), I5 =>  inp_feat(66)); 
C_38_S_5_L_5_inst : LUT6 generic map(INIT => "1101010011011100010000001101110101000001100011011100110011001100") port map( O =>C_38_S_5_L_5_out, I0 =>  inp_feat(63), I1 =>  inp_feat(51), I2 =>  inp_feat(177), I3 =>  inp_feat(482), I4 =>  inp_feat(150), I5 =>  inp_feat(64)); 
C_39_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111010111111101111100011111100111110001000100010000000") port map( O =>C_39_S_0_L_0_out, I0 =>  inp_feat(195), I1 =>  inp_feat(48), I2 =>  inp_feat(426), I3 =>  inp_feat(385), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_0_L_1_inst : LUT6 generic map(INIT => "1111001110100000111111111111111101010000000000001111111111110101") port map( O =>C_39_S_0_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(413), I2 =>  inp_feat(339), I3 =>  inp_feat(485), I4 =>  inp_feat(183), I5 =>  inp_feat(403)); 
C_39_S_0_L_2_inst : LUT6 generic map(INIT => "0111111011111000111111101100000000100000101000001000000010000000") port map( O =>C_39_S_0_L_2_out, I0 =>  inp_feat(195), I1 =>  inp_feat(232), I2 =>  inp_feat(458), I3 =>  inp_feat(482), I4 =>  inp_feat(150), I5 =>  inp_feat(463)); 
C_39_S_0_L_3_inst : LUT6 generic map(INIT => "1010100011111010111111101000000001111110000000001100000010000000") port map( O =>C_39_S_0_L_3_out, I0 =>  inp_feat(458), I1 =>  inp_feat(246), I2 =>  inp_feat(90), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_0_L_4_inst : LUT6 generic map(INIT => "0111101001110100111110101000000011101110111000000011000010000000") port map( O =>C_39_S_0_L_4_out, I0 =>  inp_feat(48), I1 =>  inp_feat(458), I2 =>  inp_feat(237), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_0_L_5_inst : LUT6 generic map(INIT => "1111110111011100110101100100100001001110101000000110100010000000") port map( O =>C_39_S_0_L_5_out, I0 =>  inp_feat(232), I1 =>  inp_feat(456), I2 =>  inp_feat(237), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_1_L_0_inst : LUT6 generic map(INIT => "1111001110100000111111111111111101110000000000001111111111110101") port map( O =>C_39_S_1_L_0_out, I0 =>  inp_feat(318), I1 =>  inp_feat(413), I2 =>  inp_feat(339), I3 =>  inp_feat(485), I4 =>  inp_feat(183), I5 =>  inp_feat(403)); 
C_39_S_1_L_1_inst : LUT6 generic map(INIT => "0100100111111010110111001010100011111110101000001100000000000000") port map( O =>C_39_S_1_L_1_out, I0 =>  inp_feat(458), I1 =>  inp_feat(456), I2 =>  inp_feat(237), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_1_L_2_inst : LUT6 generic map(INIT => "1110100011111110101010000110100000101110001110000010100000000000") port map( O =>C_39_S_1_L_2_out, I0 =>  inp_feat(124), I1 =>  inp_feat(454), I2 =>  inp_feat(432), I3 =>  inp_feat(224), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_1_L_3_inst : LUT6 generic map(INIT => "0011011001101010011010100010000011111110001010001101000010000000") port map( O =>C_39_S_1_L_3_out, I0 =>  inp_feat(458), I1 =>  inp_feat(66), I2 =>  inp_feat(237), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_1_L_4_inst : LUT6 generic map(INIT => "1111011011011100111101101100100001101110101000000110100010000000") port map( O =>C_39_S_1_L_4_out, I0 =>  inp_feat(232), I1 =>  inp_feat(456), I2 =>  inp_feat(237), I3 =>  inp_feat(482), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_39_S_1_L_5_inst : LUT6 generic map(INIT => "0010111101001110111111100000101011111110111011101101111101000010") port map( O =>C_39_S_1_L_5_out, I0 =>  inp_feat(202), I1 =>  inp_feat(332), I2 =>  inp_feat(469), I3 =>  inp_feat(115), I4 =>  inp_feat(280), I5 =>  inp_feat(20)); 
C_39_S_2_L_0_inst : LUT6 generic map(INIT => "0111111111101110111111101000000011111100000010000110100000000000") port map( O =>C_39_S_2_L_0_out, I0 =>  inp_feat(90), I1 =>  inp_feat(232), I2 =>  inp_feat(84), I3 =>  inp_feat(177), I4 =>  inp_feat(426), I5 =>  inp_feat(254)); 
C_39_S_2_L_1_inst : LUT6 generic map(INIT => "1111110011111100111111001111100000001010011011100010000010001000") port map( O =>C_39_S_2_L_1_out, I0 =>  inp_feat(232), I1 =>  inp_feat(458), I2 =>  inp_feat(482), I3 =>  inp_feat(456), I4 =>  inp_feat(426), I5 =>  inp_feat(177)); 
C_39_S_2_L_2_inst : LUT6 generic map(INIT => "1111001110001110111011101110111101110011100011100110001000101010") port map( O =>C_39_S_2_L_2_out, I0 =>  inp_feat(315), I1 =>  inp_feat(478), I2 =>  inp_feat(249), I3 =>  inp_feat(66), I4 =>  inp_feat(493), I5 =>  inp_feat(108)); 
C_39_S_2_L_3_inst : LUT6 generic map(INIT => "0001011111100010010101110000010111110111101011101111101111110111") port map( O =>C_39_S_2_L_3_out, I0 =>  inp_feat(289), I1 =>  inp_feat(149), I2 =>  inp_feat(171), I3 =>  inp_feat(482), I4 =>  inp_feat(66), I5 =>  inp_feat(183)); 
C_39_S_2_L_4_inst : LUT6 generic map(INIT => "1111111110111110111101101110000001111000111110100010100000000000") port map( O =>C_39_S_2_L_4_out, I0 =>  inp_feat(237), I1 =>  inp_feat(90), I2 =>  inp_feat(383), I3 =>  inp_feat(458), I4 =>  inp_feat(482), I5 =>  inp_feat(150)); 
C_39_S_2_L_5_inst : LUT6 generic map(INIT => "0010001000101110111111110010110111101110101111111111111100001100") port map( O =>C_39_S_2_L_5_out, I0 =>  inp_feat(475), I1 =>  inp_feat(69), I2 =>  inp_feat(426), I3 =>  inp_feat(103), I4 =>  inp_feat(124), I5 =>  inp_feat(251)); 
C_39_S_3_L_0_inst : LUT6 generic map(INIT => "1111110011110100111001001100000001010110111101101110111001000000") port map( O =>C_39_S_3_L_0_out, I0 =>  inp_feat(232), I1 =>  inp_feat(482), I2 =>  inp_feat(335), I3 =>  inp_feat(230), I4 =>  inp_feat(383), I5 =>  inp_feat(350)); 
C_39_S_3_L_1_inst : LUT6 generic map(INIT => "0101011011101010001000001110100011011110001010001100000010000000") port map( O =>C_39_S_3_L_1_out, I0 =>  inp_feat(458), I1 =>  inp_feat(456), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_3_L_2_inst : LUT6 generic map(INIT => "1011011111001010100011111110100001111110000010001100000010000000") port map( O =>C_39_S_3_L_2_out, I0 =>  inp_feat(458), I1 =>  inp_feat(456), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_3_L_3_inst : LUT6 generic map(INIT => "0011110001100010001011001110100011110110000010000000110000001000") port map( O =>C_39_S_3_L_3_out, I0 =>  inp_feat(458), I1 =>  inp_feat(232), I2 =>  inp_feat(183), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_3_L_4_inst : LUT6 generic map(INIT => "1111111101111110111110111010100001101000000010001110000010000000") port map( O =>C_39_S_3_L_4_out, I0 =>  inp_feat(232), I1 =>  inp_feat(456), I2 =>  inp_feat(245), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_3_L_5_inst : LUT6 generic map(INIT => "0011110011101100100010101110100011111110100010000110000010000000") port map( O =>C_39_S_3_L_5_out, I0 =>  inp_feat(224), I1 =>  inp_feat(458), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_4_L_0_inst : LUT6 generic map(INIT => "0111011111001110011101001110100001111110000010001010000010000000") port map( O =>C_39_S_4_L_0_out, I0 =>  inp_feat(90), I1 =>  inp_feat(458), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_4_L_1_inst : LUT6 generic map(INIT => "1011011001001010101111011110100011011110101010001100000010000000") port map( O =>C_39_S_4_L_1_out, I0 =>  inp_feat(458), I1 =>  inp_feat(456), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_4_L_2_inst : LUT6 generic map(INIT => "0111110001100100011100000110110011011110100010001010000010000000") port map( O =>C_39_S_4_L_2_out, I0 =>  inp_feat(317), I1 =>  inp_feat(458), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_4_L_3_inst : LUT6 generic map(INIT => "1100010111100100100010111110100001101110100010000110000010000000") port map( O =>C_39_S_4_L_3_out, I0 =>  inp_feat(224), I1 =>  inp_feat(458), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_4_L_4_inst : LUT6 generic map(INIT => "0101111101001100111111101010100001101000000010001110000010000000") port map( O =>C_39_S_4_L_4_out, I0 =>  inp_feat(232), I1 =>  inp_feat(456), I2 =>  inp_feat(245), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_4_L_5_inst : LUT6 generic map(INIT => "1101001110001101110101010000011110000101000011110100111101011101") port map( O =>C_39_S_4_L_5_out, I0 =>  inp_feat(69), I1 =>  inp_feat(81), I2 =>  inp_feat(139), I3 =>  inp_feat(482), I4 =>  inp_feat(150), I5 =>  inp_feat(254)); 
C_39_S_5_L_0_inst : LUT6 generic map(INIT => "1001100110000010100001011111111100000000001000101111011111111111") port map( O =>C_39_S_5_L_0_out, I0 =>  inp_feat(212), I1 =>  inp_feat(61), I2 =>  inp_feat(120), I3 =>  inp_feat(478), I4 =>  inp_feat(51), I5 =>  inp_feat(344)); 
C_39_S_5_L_1_inst : LUT6 generic map(INIT => "0000111001110111000010001101111111011111111111110100010101011111") port map( O =>C_39_S_5_L_1_out, I0 =>  inp_feat(339), I1 =>  inp_feat(492), I2 =>  inp_feat(469), I3 =>  inp_feat(378), I4 =>  inp_feat(388), I5 =>  inp_feat(404)); 
C_39_S_5_L_2_inst : LUT6 generic map(INIT => "1111111111101100101110111110100001111110110010000110000010000000") port map( O =>C_39_S_5_L_2_out, I0 =>  inp_feat(224), I1 =>  inp_feat(458), I2 =>  inp_feat(361), I3 =>  inp_feat(482), I4 =>  inp_feat(177), I5 =>  inp_feat(150)); 
C_39_S_5_L_3_inst : LUT6 generic map(INIT => "0010111111011101111111011100010000111011100011001011111101000100") port map( O =>C_39_S_5_L_3_out, I0 =>  inp_feat(100), I1 =>  inp_feat(317), I2 =>  inp_feat(232), I3 =>  inp_feat(468), I4 =>  inp_feat(176), I5 =>  inp_feat(68)); 
C_39_S_5_L_4_inst : LUT6 generic map(INIT => "1111111101001001111000110111111100001010010100101010111000001000") port map( O =>C_39_S_5_L_4_out, I0 =>  inp_feat(209), I1 =>  inp_feat(69), I2 =>  inp_feat(375), I3 =>  inp_feat(47), I4 =>  inp_feat(303), I5 =>  inp_feat(374)); 
C_39_S_5_L_5_inst : LUT6 generic map(INIT => "0011110100110011100110100010000000001000111000001101100010010000") port map( O =>C_39_S_5_L_5_out, I0 =>  inp_feat(456), I1 =>  inp_feat(483), I2 =>  inp_feat(232), I3 =>  inp_feat(482), I4 =>  inp_feat(150), I5 =>  inp_feat(254)); 
C_40_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111010111111101111100011111100111110001000100010000000") port map( O =>C_40_S_0_L_0_out, I0 =>  inp_feat(195), I1 =>  inp_feat(48), I2 =>  inp_feat(426), I3 =>  inp_feat(385), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_40_S_0_L_1_inst : LUT6 generic map(INIT => "1110011000001110000011101010111111111110111111100000111011101111") port map( O =>C_40_S_0_L_1_out, I0 =>  inp_feat(380), I1 =>  inp_feat(234), I2 =>  inp_feat(446), I3 =>  inp_feat(352), I4 =>  inp_feat(84), I5 =>  inp_feat(183)); 
C_40_S_0_L_2_inst : LUT6 generic map(INIT => "0010101001111100110111100001110100010100001101000000000011111111") port map( O =>C_40_S_0_L_2_out, I0 =>  inp_feat(454), I1 =>  inp_feat(274), I2 =>  inp_feat(0), I3 =>  inp_feat(179), I4 =>  inp_feat(317), I5 =>  inp_feat(232)); 
C_40_S_0_L_3_inst : LUT6 generic map(INIT => "1101111011111110000011101110110000000100111101000000000000000000") port map( O =>C_40_S_0_L_3_out, I0 =>  inp_feat(64), I1 =>  inp_feat(66), I2 =>  inp_feat(209), I3 =>  inp_feat(363), I4 =>  inp_feat(458), I5 =>  inp_feat(317)); 
C_40_S_0_L_4_inst : LUT6 generic map(INIT => "0111011101010001110111011111000011111111101101011101111100010011") port map( O =>C_40_S_0_L_4_out, I0 =>  inp_feat(446), I1 =>  inp_feat(152), I2 =>  inp_feat(83), I3 =>  inp_feat(218), I4 =>  inp_feat(436), I5 =>  inp_feat(503)); 
C_40_S_0_L_5_inst : LUT6 generic map(INIT => "1101100011111111110111011111100001111000111100000010100010100000") port map( O =>C_40_S_0_L_5_out, I0 =>  inp_feat(89), I1 =>  inp_feat(67), I2 =>  inp_feat(509), I3 =>  inp_feat(94), I4 =>  inp_feat(504), I5 =>  inp_feat(335)); 
C_40_S_1_L_0_inst : LUT6 generic map(INIT => "1110011000001110000011101010111111111110111111100000111011101111") port map( O =>C_40_S_1_L_0_out, I0 =>  inp_feat(380), I1 =>  inp_feat(234), I2 =>  inp_feat(446), I3 =>  inp_feat(352), I4 =>  inp_feat(84), I5 =>  inp_feat(183)); 
C_40_S_1_L_1_inst : LUT6 generic map(INIT => "0010101001111100110111100001110100010100001101000000000011111111") port map( O =>C_40_S_1_L_1_out, I0 =>  inp_feat(454), I1 =>  inp_feat(274), I2 =>  inp_feat(0), I3 =>  inp_feat(179), I4 =>  inp_feat(317), I5 =>  inp_feat(232)); 
C_40_S_1_L_2_inst : LUT6 generic map(INIT => "1101111011111110000011101110110000000100111101000000000000000000") port map( O =>C_40_S_1_L_2_out, I0 =>  inp_feat(64), I1 =>  inp_feat(66), I2 =>  inp_feat(209), I3 =>  inp_feat(363), I4 =>  inp_feat(458), I5 =>  inp_feat(317)); 
C_40_S_1_L_3_inst : LUT6 generic map(INIT => "0111011101010001110111011111000011111111101101011101111100010011") port map( O =>C_40_S_1_L_3_out, I0 =>  inp_feat(446), I1 =>  inp_feat(152), I2 =>  inp_feat(83), I3 =>  inp_feat(218), I4 =>  inp_feat(436), I5 =>  inp_feat(503)); 
C_40_S_1_L_4_inst : LUT6 generic map(INIT => "1101100011111111110111011111100001111000111100000010100010100000") port map( O =>C_40_S_1_L_4_out, I0 =>  inp_feat(89), I1 =>  inp_feat(67), I2 =>  inp_feat(509), I3 =>  inp_feat(94), I4 =>  inp_feat(504), I5 =>  inp_feat(335)); 
C_40_S_1_L_5_inst : LUT6 generic map(INIT => "0101101111111110010010001111100000000010111110001000000000000000") port map( O =>C_40_S_1_L_5_out, I0 =>  inp_feat(150), I1 =>  inp_feat(232), I2 =>  inp_feat(458), I3 =>  inp_feat(37), I4 =>  inp_feat(315), I5 =>  inp_feat(81)); 
C_40_S_2_L_0_inst : LUT6 generic map(INIT => "0110110111111011111001111101001101111101111111000000001010110010") port map( O =>C_40_S_2_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(432), I2 =>  inp_feat(195), I3 =>  inp_feat(147), I4 =>  inp_feat(482), I5 =>  inp_feat(90)); 
C_40_S_2_L_1_inst : LUT6 generic map(INIT => "1010000110101101011110111001110101010011111111110000000011100000") port map( O =>C_40_S_2_L_1_out, I0 =>  inp_feat(48), I1 =>  inp_feat(289), I2 =>  inp_feat(448), I3 =>  inp_feat(147), I4 =>  inp_feat(482), I5 =>  inp_feat(90)); 
C_40_S_2_L_2_inst : LUT6 generic map(INIT => "0011001100100011000001000111001111111110101111100100111011111110") port map( O =>C_40_S_2_L_2_out, I0 =>  inp_feat(385), I1 =>  inp_feat(151), I2 =>  inp_feat(242), I3 =>  inp_feat(15), I4 =>  inp_feat(4), I5 =>  inp_feat(33)); 
C_40_S_2_L_3_inst : LUT6 generic map(INIT => "1101110111101111101011000000110001100110011001010000101000000000") port map( O =>C_40_S_2_L_3_out, I0 =>  inp_feat(492), I1 =>  inp_feat(17), I2 =>  inp_feat(244), I3 =>  inp_feat(177), I4 =>  inp_feat(315), I5 =>  inp_feat(81)); 
C_40_S_2_L_4_inst : LUT6 generic map(INIT => "0100001000011011000001101000100111111111011011000000111011111010") port map( O =>C_40_S_2_L_4_out, I0 =>  inp_feat(145), I1 =>  inp_feat(239), I2 =>  inp_feat(4), I3 =>  inp_feat(334), I4 =>  inp_feat(218), I5 =>  inp_feat(479)); 
C_40_S_2_L_5_inst : LUT6 generic map(INIT => "1110111010100000011111101010000000011001000010001111111110000000") port map( O =>C_40_S_2_L_5_out, I0 =>  inp_feat(346), I1 =>  inp_feat(426), I2 =>  inp_feat(473), I3 =>  inp_feat(458), I4 =>  inp_feat(88), I5 =>  inp_feat(0)); 
C_40_S_3_L_0_inst : LUT6 generic map(INIT => "0000011001101101000000110011111111101111011111110110111101011111") port map( O =>C_40_S_3_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(16), I2 =>  inp_feat(253), I3 =>  inp_feat(4), I4 =>  inp_feat(105), I5 =>  inp_feat(33)); 
C_40_S_3_L_1_inst : LUT6 generic map(INIT => "0101101111111111001100110011110111111110111111001111100001101000") port map( O =>C_40_S_3_L_1_out, I0 =>  inp_feat(510), I1 =>  inp_feat(92), I2 =>  inp_feat(382), I3 =>  inp_feat(435), I4 =>  inp_feat(130), I5 =>  inp_feat(419)); 
C_40_S_3_L_2_inst : LUT6 generic map(INIT => "1110011110101110100001111111111110100101110111110010001100000010") port map( O =>C_40_S_3_L_2_out, I0 =>  inp_feat(90), I1 =>  inp_feat(157), I2 =>  inp_feat(126), I3 =>  inp_feat(95), I4 =>  inp_feat(383), I5 =>  inp_feat(230)); 
C_40_S_3_L_3_inst : LUT6 generic map(INIT => "0100110000111111010001110110111111111100111010111111111001001010") port map( O =>C_40_S_3_L_3_out, I0 =>  inp_feat(445), I1 =>  inp_feat(493), I2 =>  inp_feat(407), I3 =>  inp_feat(75), I4 =>  inp_feat(162), I5 =>  inp_feat(479)); 
C_40_S_3_L_4_inst : LUT6 generic map(INIT => "1111111011100100110110001110000000001100101010001110000011001000") port map( O =>C_40_S_3_L_4_out, I0 =>  inp_feat(150), I1 =>  inp_feat(237), I2 =>  inp_feat(232), I3 =>  inp_feat(447), I4 =>  inp_feat(54), I5 =>  inp_feat(413)); 
C_40_S_3_L_5_inst : LUT6 generic map(INIT => "0011101000110010101010011111100011111111111110000011011011111010") port map( O =>C_40_S_3_L_5_out, I0 =>  inp_feat(470), I1 =>  inp_feat(422), I2 =>  inp_feat(371), I3 =>  inp_feat(500), I4 =>  inp_feat(231), I5 =>  inp_feat(111)); 
C_40_S_4_L_0_inst : LUT6 generic map(INIT => "1111000011101010111011101110110010100010001100111110111111100110") port map( O =>C_40_S_4_L_0_out, I0 =>  inp_feat(203), I1 =>  inp_feat(418), I2 =>  inp_feat(345), I3 =>  inp_feat(489), I4 =>  inp_feat(220), I5 =>  inp_feat(290)); 
C_40_S_4_L_1_inst : LUT6 generic map(INIT => "1111111100001010111000101000100000100000011011001100010000000000") port map( O =>C_40_S_4_L_1_out, I0 =>  inp_feat(482), I1 =>  inp_feat(150), I2 =>  inp_feat(398), I3 =>  inp_feat(237), I4 =>  inp_feat(66), I5 =>  inp_feat(245)); 
C_40_S_4_L_2_inst : LUT6 generic map(INIT => "0111011101101101000011101110100010101110001010000000000010000000") port map( O =>C_40_S_4_L_2_out, I0 =>  inp_feat(232), I1 =>  inp_feat(456), I2 =>  inp_feat(463), I3 =>  inp_feat(45), I4 =>  inp_feat(230), I5 =>  inp_feat(383)); 
C_40_S_4_L_3_inst : LUT6 generic map(INIT => "1111111101010101000010100011111100110111110101110010000010111010") port map( O =>C_40_S_4_L_3_out, I0 =>  inp_feat(64), I1 =>  inp_feat(454), I2 =>  inp_feat(339), I3 =>  inp_feat(204), I4 =>  inp_feat(66), I5 =>  inp_feat(7)); 
C_40_S_4_L_4_inst : LUT6 generic map(INIT => "0101001010100010011101100000111011111111011011101110000000000000") port map( O =>C_40_S_4_L_4_out, I0 =>  inp_feat(232), I1 =>  inp_feat(84), I2 =>  inp_feat(31), I3 =>  inp_feat(335), I4 =>  inp_feat(137), I5 =>  inp_feat(344)); 
C_40_S_4_L_5_inst : LUT6 generic map(INIT => "0101101111100010110100100111111011011011111111001010101011100000") port map( O =>C_40_S_4_L_5_out, I0 =>  inp_feat(445), I1 =>  inp_feat(334), I2 =>  inp_feat(391), I3 =>  inp_feat(83), I4 =>  inp_feat(207), I5 =>  inp_feat(220)); 
C_40_S_5_L_0_inst : LUT6 generic map(INIT => "1101101110100011111100110111111101110111111110111111111111110010") port map( O =>C_40_S_5_L_0_out, I0 =>  inp_feat(179), I1 =>  inp_feat(86), I2 =>  inp_feat(391), I3 =>  inp_feat(83), I4 =>  inp_feat(207), I5 =>  inp_feat(220)); 
C_40_S_5_L_1_inst : LUT6 generic map(INIT => "1010001110010010111110110000000001001110111100101101000000000000") port map( O =>C_40_S_5_L_1_out, I0 =>  inp_feat(357), I1 =>  inp_feat(313), I2 =>  inp_feat(315), I3 =>  inp_feat(232), I4 =>  inp_feat(66), I5 =>  inp_feat(245)); 
C_40_S_5_L_2_inst : LUT6 generic map(INIT => "1111100010101100101110101010111000010011111111010000110001000000") port map( O =>C_40_S_5_L_2_out, I0 =>  inp_feat(90), I1 =>  inp_feat(357), I2 =>  inp_feat(312), I3 =>  inp_feat(315), I4 =>  inp_feat(50), I5 =>  inp_feat(244)); 
C_40_S_5_L_3_inst : LUT6 generic map(INIT => "0001010110010100010100011100010100010001110100111111010100010100") port map( O =>C_40_S_5_L_3_out, I0 =>  inp_feat(52), I1 =>  inp_feat(224), I2 =>  inp_feat(290), I3 =>  inp_feat(242), I4 =>  inp_feat(78), I5 =>  inp_feat(109)); 
C_40_S_5_L_4_inst : LUT6 generic map(INIT => "0111000000001100111110000000010011101111111011101110100000101100") port map( O =>C_40_S_5_L_4_out, I0 =>  inp_feat(237), I1 =>  inp_feat(458), I2 =>  inp_feat(473), I3 =>  inp_feat(230), I4 =>  inp_feat(65), I5 =>  inp_feat(303)); 
C_40_S_5_L_5_inst : LUT6 generic map(INIT => "1111010111101111001101111111111100001001110011011111011111111111") port map( O =>C_40_S_5_L_5_out, I0 =>  inp_feat(395), I1 =>  inp_feat(510), I2 =>  inp_feat(394), I3 =>  inp_feat(179), I4 =>  inp_feat(419), I5 =>  inp_feat(231)); 
C_41_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111110111111101110100011111110111110001100100010000000") port map( O =>C_41_S_0_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(48), I2 =>  inp_feat(426), I3 =>  inp_feat(385), I4 =>  inp_feat(383), I5 =>  inp_feat(150)); 
C_41_S_0_L_1_inst : LUT6 generic map(INIT => "1000110011000000000101000110000011111011110111101110100000000000") port map( O =>C_41_S_0_L_1_out, I0 =>  inp_feat(84), I1 =>  inp_feat(232), I2 =>  inp_feat(473), I3 =>  inp_feat(66), I4 =>  inp_feat(383), I5 =>  inp_feat(46)); 
C_41_S_0_L_2_inst : LUT6 generic map(INIT => "0101011111100111110001001110011111011111111111001111111011001000") port map( O =>C_41_S_0_L_2_out, I0 =>  inp_feat(296), I1 =>  inp_feat(105), I2 =>  inp_feat(164), I3 =>  inp_feat(338), I4 =>  inp_feat(183), I5 =>  inp_feat(46)); 
C_41_S_0_L_3_inst : LUT6 generic map(INIT => "1101110111010100111101001111011111111101110011111111111101011101") port map( O =>C_41_S_0_L_3_out, I0 =>  inp_feat(277), I1 =>  inp_feat(286), I2 =>  inp_feat(232), I3 =>  inp_feat(296), I4 =>  inp_feat(246), I5 =>  inp_feat(275)); 
C_41_S_0_L_4_inst : LUT6 generic map(INIT => "0100010111100000110001001111011110101100111110001111000011111000") port map( O =>C_41_S_0_L_4_out, I0 =>  inp_feat(166), I1 =>  inp_feat(341), I2 =>  inp_feat(485), I3 =>  inp_feat(277), I4 =>  inp_feat(187), I5 =>  inp_feat(275)); 
C_41_S_0_L_5_inst : LUT6 generic map(INIT => "1100111011001110111101111000111101011101001010101000111100000000") port map( O =>C_41_S_0_L_5_out, I0 =>  inp_feat(90), I1 =>  inp_feat(445), I2 =>  inp_feat(115), I3 =>  inp_feat(66), I4 =>  inp_feat(237), I5 =>  inp_feat(492)); 
C_41_S_1_L_0_inst : LUT6 generic map(INIT => "1000110011000000000101000110000011111011110111101110100000000000") port map( O =>C_41_S_1_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(232), I2 =>  inp_feat(473), I3 =>  inp_feat(66), I4 =>  inp_feat(383), I5 =>  inp_feat(46)); 
C_41_S_1_L_1_inst : LUT6 generic map(INIT => "0101011111100111110001001110011111011111111111001111111011001000") port map( O =>C_41_S_1_L_1_out, I0 =>  inp_feat(296), I1 =>  inp_feat(105), I2 =>  inp_feat(164), I3 =>  inp_feat(338), I4 =>  inp_feat(183), I5 =>  inp_feat(46)); 
C_41_S_1_L_2_inst : LUT6 generic map(INIT => "1101110111010100111101001111011111111101110011111111111101011101") port map( O =>C_41_S_1_L_2_out, I0 =>  inp_feat(277), I1 =>  inp_feat(286), I2 =>  inp_feat(232), I3 =>  inp_feat(296), I4 =>  inp_feat(246), I5 =>  inp_feat(275)); 
C_41_S_1_L_3_inst : LUT6 generic map(INIT => "0100010111100000110001001111011110101100111110001111000011111000") port map( O =>C_41_S_1_L_3_out, I0 =>  inp_feat(166), I1 =>  inp_feat(341), I2 =>  inp_feat(485), I3 =>  inp_feat(277), I4 =>  inp_feat(187), I5 =>  inp_feat(275)); 
C_41_S_1_L_4_inst : LUT6 generic map(INIT => "1100111011001110111101111000111101011101001010101000111100000000") port map( O =>C_41_S_1_L_4_out, I0 =>  inp_feat(90), I1 =>  inp_feat(445), I2 =>  inp_feat(115), I3 =>  inp_feat(66), I4 =>  inp_feat(237), I5 =>  inp_feat(492)); 
C_41_S_1_L_5_inst : LUT6 generic map(INIT => "0100111101111010010101100000101011111111111111101111111001001011") port map( O =>C_41_S_1_L_5_out, I0 =>  inp_feat(277), I1 =>  inp_feat(44), I2 =>  inp_feat(270), I3 =>  inp_feat(173), I4 =>  inp_feat(180), I5 =>  inp_feat(389)); 
C_41_S_2_L_0_inst : LUT6 generic map(INIT => "1111110101111111101111011111110001011111001101110101101011110000") port map( O =>C_41_S_2_L_0_out, I0 =>  inp_feat(189), I1 =>  inp_feat(217), I2 =>  inp_feat(387), I3 =>  inp_feat(116), I4 =>  inp_feat(473), I5 =>  inp_feat(232)); 
C_41_S_2_L_1_inst : LUT6 generic map(INIT => "1011110010101101100000001111001000101110001011101000000011110001") port map( O =>C_41_S_2_L_1_out, I0 =>  inp_feat(492), I1 =>  inp_feat(17), I2 =>  inp_feat(426), I3 =>  inp_feat(338), I4 =>  inp_feat(177), I5 =>  inp_feat(383)); 
C_41_S_2_L_2_inst : LUT6 generic map(INIT => "0001100001100110110101010111011010000010111010101111110011101000") port map( O =>C_41_S_2_L_2_out, I0 =>  inp_feat(150), I1 =>  inp_feat(64), I2 =>  inp_feat(385), I3 =>  inp_feat(164), I4 =>  inp_feat(183), I5 =>  inp_feat(46)); 
C_41_S_2_L_3_inst : LUT6 generic map(INIT => "0011001111110010111110111011011111101011111101101111111111111111") port map( O =>C_41_S_2_L_3_out, I0 =>  inp_feat(23), I1 =>  inp_feat(124), I2 =>  inp_feat(310), I3 =>  inp_feat(166), I4 =>  inp_feat(387), I5 =>  inp_feat(320)); 
C_41_S_2_L_4_inst : LUT6 generic map(INIT => "1010101011101100100111100101100011111100111100001111110000000000") port map( O =>C_41_S_2_L_4_out, I0 =>  inp_feat(1), I1 =>  inp_feat(159), I2 =>  inp_feat(163), I3 =>  inp_feat(237), I4 =>  inp_feat(344), I5 =>  inp_feat(218)); 
C_41_S_2_L_5_inst : LUT6 generic map(INIT => "1110111111101110101011111101111101000000110111111111111110001111") port map( O =>C_41_S_2_L_5_out, I0 =>  inp_feat(66), I1 =>  inp_feat(232), I2 =>  inp_feat(465), I3 =>  inp_feat(129), I4 =>  inp_feat(410), I5 =>  inp_feat(286)); 
C_41_S_3_L_0_inst : LUT6 generic map(INIT => "1001111001101100000000000111010001011000011010000000000010100000") port map( O =>C_41_S_3_L_0_out, I0 =>  inp_feat(482), I1 =>  inp_feat(237), I2 =>  inp_feat(150), I3 =>  inp_feat(93), I4 =>  inp_feat(137), I5 =>  inp_feat(383)); 
C_41_S_3_L_1_inst : LUT6 generic map(INIT => "0001110010000001001001111111010011111111101011011001111010110101") port map( O =>C_41_S_3_L_1_out, I0 =>  inp_feat(453), I1 =>  inp_feat(195), I2 =>  inp_feat(245), I3 =>  inp_feat(398), I4 =>  inp_feat(407), I5 =>  inp_feat(20)); 
C_41_S_3_L_2_inst : LUT6 generic map(INIT => "1110100101111100100110101111111100011111101111100010000111111111") port map( O =>C_41_S_3_L_2_out, I0 =>  inp_feat(317), I1 =>  inp_feat(253), I2 =>  inp_feat(494), I3 =>  inp_feat(325), I4 =>  inp_feat(361), I5 =>  inp_feat(176)); 
C_41_S_3_L_3_inst : LUT6 generic map(INIT => "1101111010001011110111111100111101001110011011111111111111001111") port map( O =>C_41_S_3_L_3_out, I0 =>  inp_feat(306), I1 =>  inp_feat(91), I2 =>  inp_feat(107), I3 =>  inp_feat(164), I4 =>  inp_feat(25), I5 =>  inp_feat(113)); 
C_41_S_3_L_4_inst : LUT6 generic map(INIT => "0000010100000100101011010010110111011111001101011111111101011110") port map( O =>C_41_S_3_L_4_out, I0 =>  inp_feat(368), I1 =>  inp_feat(200), I2 =>  inp_feat(115), I3 =>  inp_feat(445), I4 =>  inp_feat(77), I5 =>  inp_feat(221)); 
C_41_S_3_L_5_inst : LUT6 generic map(INIT => "1010011010001100101011111111001011101011111010001111111010000000") port map( O =>C_41_S_3_L_5_out, I0 =>  inp_feat(214), I1 =>  inp_feat(42), I2 =>  inp_feat(352), I3 =>  inp_feat(4), I4 =>  inp_feat(14), I5 =>  inp_feat(389)); 
C_41_S_4_L_0_inst : LUT6 generic map(INIT => "1110001111101110011001111010101111111111111110111111101110100010") port map( O =>C_41_S_4_L_0_out, I0 =>  inp_feat(266), I1 =>  inp_feat(427), I2 =>  inp_feat(75), I3 =>  inp_feat(180), I4 =>  inp_feat(91), I5 =>  inp_feat(141)); 
C_41_S_4_L_1_inst : LUT6 generic map(INIT => "1110011100111111110000001111110011100000110111101000000010100000") port map( O =>C_41_S_4_L_1_out, I0 =>  inp_feat(257), I1 =>  inp_feat(315), I2 =>  inp_feat(84), I3 =>  inp_feat(183), I4 =>  inp_feat(468), I5 =>  inp_feat(335)); 
C_41_S_4_L_2_inst : LUT6 generic map(INIT => "1100111110101100101011101101110000101010001011001111110011111000") port map( O =>C_41_S_4_L_2_out, I0 =>  inp_feat(176), I1 =>  inp_feat(383), I2 =>  inp_feat(129), I3 =>  inp_feat(295), I4 =>  inp_feat(410), I5 =>  inp_feat(286)); 
C_41_S_4_L_3_inst : LUT6 generic map(INIT => "0010010000001111110011000010100010110100101000101111100010100000") port map( O =>C_41_S_4_L_3_out, I0 =>  inp_feat(482), I1 =>  inp_feat(237), I2 =>  inp_feat(200), I3 =>  inp_feat(4), I4 =>  inp_feat(14), I5 =>  inp_feat(503)); 
C_41_S_4_L_4_inst : LUT6 generic map(INIT => "1110001011110011101010001010101010110000100000010010000110000000") port map( O =>C_41_S_4_L_4_out, I0 =>  inp_feat(317), I1 =>  inp_feat(251), I2 =>  inp_feat(430), I3 =>  inp_feat(107), I4 =>  inp_feat(468), I5 =>  inp_feat(398)); 
C_41_S_4_L_5_inst : LUT6 generic map(INIT => "1110101001101000100111101110110001010101011110101111101010100000") port map( O =>C_41_S_4_L_5_out, I0 =>  inp_feat(264), I1 =>  inp_feat(176), I2 =>  inp_feat(383), I3 =>  inp_feat(363), I4 =>  inp_feat(410), I5 =>  inp_feat(429)); 
C_41_S_5_L_0_inst : LUT6 generic map(INIT => "0110010001111110100011001000110011100110001011000000000110000100") port map( O =>C_41_S_5_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(232), I2 =>  inp_feat(278), I3 =>  inp_feat(413), I4 =>  inp_feat(42), I5 =>  inp_feat(286)); 
C_41_S_5_L_1_inst : LUT6 generic map(INIT => "0111100111101110100100001110101011101101111101100000100010001010") port map( O =>C_41_S_5_L_1_out, I0 =>  inp_feat(442), I1 =>  inp_feat(454), I2 =>  inp_feat(510), I3 =>  inp_feat(269), I4 =>  inp_feat(55), I5 =>  inp_feat(332)); 
C_41_S_5_L_2_inst : LUT6 generic map(INIT => "1100111111101110111011111110111100011100011010101011111111111111") port map( O =>C_41_S_5_L_2_out, I0 =>  inp_feat(89), I1 =>  inp_feat(378), I2 =>  inp_feat(289), I3 =>  inp_feat(244), I4 =>  inp_feat(320), I5 =>  inp_feat(111)); 
C_41_S_5_L_3_inst : LUT6 generic map(INIT => "1100100001011000111100100001100000101100110111011110110011000000") port map( O =>C_41_S_5_L_3_out, I0 =>  inp_feat(150), I1 =>  inp_feat(315), I2 =>  inp_feat(386), I3 =>  inp_feat(375), I4 =>  inp_feat(349), I5 =>  inp_feat(180)); 
C_41_S_5_L_4_inst : LUT6 generic map(INIT => "0011101010001111011001011111111100110111011000101011000111101111") port map( O =>C_41_S_5_L_4_out, I0 =>  inp_feat(180), I1 =>  inp_feat(141), I2 =>  inp_feat(339), I3 =>  inp_feat(101), I4 =>  inp_feat(83), I5 =>  inp_feat(113)); 
C_41_S_5_L_5_inst : LUT6 generic map(INIT => "1101111101011111101111111111111101101110111111110011111111111110") port map( O =>C_41_S_5_L_5_out, I0 =>  inp_feat(105), I1 =>  inp_feat(335), I2 =>  inp_feat(288), I3 =>  inp_feat(140), I4 =>  inp_feat(94), I5 =>  inp_feat(472)); 
C_42_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000") port map( O =>C_42_S_0_L_0_out, I0 =>  inp_feat(453), I1 =>  inp_feat(234), I2 =>  inp_feat(306), I3 =>  inp_feat(10), I4 =>  inp_feat(182), I5 =>  inp_feat(285)); 
C_42_S_0_L_1_inst : LUT6 generic map(INIT => "1010101110011000000011110000000000000000010110000000011100000100") port map( O =>C_42_S_0_L_1_out, I0 =>  inp_feat(91), I1 =>  inp_feat(320), I2 =>  inp_feat(190), I3 =>  inp_feat(10), I4 =>  inp_feat(399), I5 =>  inp_feat(194)); 
C_42_S_0_L_2_inst : LUT6 generic map(INIT => "0100011001111110011101110110111111101110111111110111111111101111") port map( O =>C_42_S_0_L_2_out, I0 =>  inp_feat(453), I1 =>  inp_feat(123), I2 =>  inp_feat(317), I3 =>  inp_feat(74), I4 =>  inp_feat(476), I5 =>  inp_feat(147)); 
C_42_S_0_L_3_inst : LUT6 generic map(INIT => "1110111011111100101001100010110000001110010111100010110000000000") port map( O =>C_42_S_0_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(395), I2 =>  inp_feat(324), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(369)); 
C_42_S_0_L_4_inst : LUT6 generic map(INIT => "0000000000010111011011111110111101111010001010111111111111111111") port map( O =>C_42_S_0_L_4_out, I0 =>  inp_feat(511), I1 =>  inp_feat(65), I2 =>  inp_feat(13), I3 =>  inp_feat(74), I4 =>  inp_feat(476), I5 =>  inp_feat(469)); 
C_42_S_0_L_5_inst : LUT6 generic map(INIT => "0111111111110010111111101010100011111111111111001110010000000000") port map( O =>C_42_S_0_L_5_out, I0 =>  inp_feat(234), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_1_L_0_inst : LUT6 generic map(INIT => "0101101011111101010101111111111111111110111111011111111111111111") port map( O =>C_42_S_1_L_0_out, I0 =>  inp_feat(246), I1 =>  inp_feat(83), I2 =>  inp_feat(74), I3 =>  inp_feat(50), I4 =>  inp_feat(378), I5 =>  inp_feat(451)); 
C_42_S_1_L_1_inst : LUT6 generic map(INIT => "1111111011101100111111001000100001100110010001001000000010001000") port map( O =>C_42_S_1_L_1_out, I0 =>  inp_feat(91), I1 =>  inp_feat(20), I2 =>  inp_feat(488), I3 =>  inp_feat(10), I4 =>  inp_feat(285), I5 =>  inp_feat(30)); 
C_42_S_1_L_2_inst : LUT6 generic map(INIT => "0101100111111110111111001010100001100010111110101000000000000000") port map( O =>C_42_S_1_L_2_out, I0 =>  inp_feat(494), I1 =>  inp_feat(123), I2 =>  inp_feat(207), I3 =>  inp_feat(507), I4 =>  inp_feat(234), I5 =>  inp_feat(225)); 
C_42_S_1_L_3_inst : LUT6 generic map(INIT => "1000110101000011110011001101100011011001110110011101000011110100") port map( O =>C_42_S_1_L_3_out, I0 =>  inp_feat(228), I1 =>  inp_feat(1), I2 =>  inp_feat(410), I3 =>  inp_feat(74), I4 =>  inp_feat(84), I5 =>  inp_feat(469)); 
C_42_S_1_L_4_inst : LUT6 generic map(INIT => "0110010100001100000001011110111111111111111111011101111111011111") port map( O =>C_42_S_1_L_4_out, I0 =>  inp_feat(51), I1 =>  inp_feat(374), I2 =>  inp_feat(317), I3 =>  inp_feat(74), I4 =>  inp_feat(476), I5 =>  inp_feat(147)); 
C_42_S_1_L_5_inst : LUT6 generic map(INIT => "1011110111110100101110110011101100001010011100100010101000000010") port map( O =>C_42_S_1_L_5_out, I0 =>  inp_feat(136), I1 =>  inp_feat(143), I2 =>  inp_feat(365), I3 =>  inp_feat(285), I4 =>  inp_feat(179), I5 =>  inp_feat(17)); 
C_42_S_2_L_0_inst : LUT6 generic map(INIT => "0100011100101111000101011110111111101111111011110101111111111111") port map( O =>C_42_S_2_L_0_out, I0 =>  inp_feat(289), I1 =>  inp_feat(273), I2 =>  inp_feat(317), I3 =>  inp_feat(74), I4 =>  inp_feat(476), I5 =>  inp_feat(147)); 
C_42_S_2_L_1_inst : LUT6 generic map(INIT => "1111111110111001111101011101010011111111111110001100010000000000") port map( O =>C_42_S_2_L_1_out, I0 =>  inp_feat(385), I1 =>  inp_feat(285), I2 =>  inp_feat(494), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_2_L_2_inst : LUT6 generic map(INIT => "0010001100100000011001111010001010010001111010001011000110101000") port map( O =>C_42_S_2_L_2_out, I0 =>  inp_feat(510), I1 =>  inp_feat(431), I2 =>  inp_feat(279), I3 =>  inp_feat(391), I4 =>  inp_feat(84), I5 =>  inp_feat(469)); 
C_42_S_2_L_3_inst : LUT6 generic map(INIT => "1111111111110100111111110101010100000000000000001111111010000000") port map( O =>C_42_S_2_L_3_out, I0 =>  inp_feat(307), I1 =>  inp_feat(21), I2 =>  inp_feat(480), I3 =>  inp_feat(10), I4 =>  inp_feat(1), I5 =>  inp_feat(194)); 
C_42_S_2_L_4_inst : LUT6 generic map(INIT => "0000000100100110111010110000001011111111111110110001111100000000") port map( O =>C_42_S_2_L_4_out, I0 =>  inp_feat(485), I1 =>  inp_feat(338), I2 =>  inp_feat(130), I3 =>  inp_feat(21), I4 =>  inp_feat(494), I5 =>  inp_feat(24)); 
C_42_S_2_L_5_inst : LUT6 generic map(INIT => "0111111101111111011101110100111011101100001111101000000010000000") port map( O =>C_42_S_2_L_5_out, I0 =>  inp_feat(91), I1 =>  inp_feat(10), I2 =>  inp_feat(503), I3 =>  inp_feat(374), I4 =>  inp_feat(21), I5 =>  inp_feat(494)); 
C_42_S_3_L_0_inst : LUT6 generic map(INIT => "0010100110001000101011001000110011111100111010101110110011111110") port map( O =>C_42_S_3_L_0_out, I0 =>  inp_feat(0), I1 =>  inp_feat(207), I2 =>  inp_feat(75), I3 =>  inp_feat(74), I4 =>  inp_feat(249), I5 =>  inp_feat(81)); 
C_42_S_3_L_1_inst : LUT6 generic map(INIT => "1110110110011011100111111010101111111101111100011000001100000010") port map( O =>C_42_S_3_L_1_out, I0 =>  inp_feat(182), I1 =>  inp_feat(287), I2 =>  inp_feat(20), I3 =>  inp_feat(234), I4 =>  inp_feat(10), I5 =>  inp_feat(285)); 
C_42_S_3_L_2_inst : LUT6 generic map(INIT => "0000010100110101010111010001110111010111111111111100111110111111") port map( O =>C_42_S_3_L_2_out, I0 =>  inp_feat(199), I1 =>  inp_feat(76), I2 =>  inp_feat(74), I3 =>  inp_feat(391), I4 =>  inp_feat(470), I5 =>  inp_feat(451)); 
C_42_S_3_L_3_inst : LUT6 generic map(INIT => "1111111111001100111111011101010111000100010011111010000000000000") port map( O =>C_42_S_3_L_3_out, I0 =>  inp_feat(363), I1 =>  inp_feat(182), I2 =>  inp_feat(123), I3 =>  inp_feat(494), I4 =>  inp_feat(371), I5 =>  inp_feat(186)); 
C_42_S_3_L_4_inst : LUT6 generic map(INIT => "0110011111000100101011010010001001010101110001001010110110100000") port map( O =>C_42_S_3_L_4_out, I0 =>  inp_feat(98), I1 =>  inp_feat(183), I2 =>  inp_feat(493), I3 =>  inp_feat(312), I4 =>  inp_feat(306), I5 =>  inp_feat(404)); 
C_42_S_3_L_5_inst : LUT6 generic map(INIT => "1100001010100110100010110000001000000000000001000001111000000000") port map( O =>C_42_S_3_L_5_out, I0 =>  inp_feat(272), I1 =>  inp_feat(131), I2 =>  inp_feat(448), I3 =>  inp_feat(182), I4 =>  inp_feat(499), I5 =>  inp_feat(467)); 
C_42_S_4_L_0_inst : LUT6 generic map(INIT => "1101101100011011101111110011010111011011000011011101001100000000") port map( O =>C_42_S_4_L_0_out, I0 =>  inp_feat(476), I1 =>  inp_feat(50), I2 =>  inp_feat(123), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_4_L_1_inst : LUT6 generic map(INIT => "0001010111010010111111101010100011011111111111001110010000000000") port map( O =>C_42_S_4_L_1_out, I0 =>  inp_feat(234), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_4_L_2_inst : LUT6 generic map(INIT => "0001111001110110000101101011100000111110111111111001110011101111") port map( O =>C_42_S_4_L_2_out, I0 =>  inp_feat(227), I1 =>  inp_feat(47), I2 =>  inp_feat(48), I3 =>  inp_feat(447), I4 =>  inp_feat(391), I5 =>  inp_feat(246)); 
C_42_S_4_L_3_inst : LUT6 generic map(INIT => "1111111101100110011101001000000011111111101010001110010000000000") port map( O =>C_42_S_4_L_3_out, I0 =>  inp_feat(10), I1 =>  inp_feat(285), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_4_L_4_inst : LUT6 generic map(INIT => "0000100011110001101110111101000011011011110101011000000000000000") port map( O =>C_42_S_4_L_4_out, I0 =>  inp_feat(248), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_4_L_5_inst : LUT6 generic map(INIT => "1001010111111010011101101010100010010110011111101110010000000000") port map( O =>C_42_S_4_L_5_out, I0 =>  inp_feat(234), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_5_L_0_inst : LUT6 generic map(INIT => "0100111110001001110111101011000011111101010100011000000000000000") port map( O =>C_42_S_5_L_0_out, I0 =>  inp_feat(123), I1 =>  inp_feat(248), I2 =>  inp_feat(285), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_5_L_1_inst : LUT6 generic map(INIT => "0111111111111010011101101010100011110110111111101110010000000000") port map( O =>C_42_S_5_L_1_out, I0 =>  inp_feat(234), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_5_L_2_inst : LUT6 generic map(INIT => "1010110011110001110110011101000011011011110101011000000000000000") port map( O =>C_42_S_5_L_2_out, I0 =>  inp_feat(248), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_5_L_3_inst : LUT6 generic map(INIT => "1001101101100110011101101000000001111111001010001110010000000000") port map( O =>C_42_S_5_L_3_out, I0 =>  inp_feat(10), I1 =>  inp_feat(285), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_5_L_4_inst : LUT6 generic map(INIT => "0111101101010111100011110011010101011011000001011101001100000000") port map( O =>C_42_S_5_L_4_out, I0 =>  inp_feat(476), I1 =>  inp_feat(50), I2 =>  inp_feat(123), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_42_S_5_L_5_inst : LUT6 generic map(INIT => "1100110110110101011100111101000011111111101101011000000000000000") port map( O =>C_42_S_5_L_5_out, I0 =>  inp_feat(248), I1 =>  inp_feat(507), I2 =>  inp_feat(292), I3 =>  inp_feat(182), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_43_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111111110100011111110111010001110110010000000") port map( O =>C_43_S_0_L_0_out, I0 =>  inp_feat(91), I1 =>  inp_feat(234), I2 =>  inp_feat(306), I3 =>  inp_feat(10), I4 =>  inp_feat(182), I5 =>  inp_feat(285)); 
C_43_S_0_L_1_inst : LUT6 generic map(INIT => "1111111010111111111111101110000000100000001111001110100010000000") port map( O =>C_43_S_0_L_1_out, I0 =>  inp_feat(120), I1 =>  inp_feat(381), I2 =>  inp_feat(210), I3 =>  inp_feat(487), I4 =>  inp_feat(434), I5 =>  inp_feat(91)); 
C_43_S_0_L_2_inst : LUT6 generic map(INIT => "0000110111011101111101111101010011111111110111101111110000001100") port map( O =>C_43_S_0_L_2_out, I0 =>  inp_feat(228), I1 =>  inp_feat(470), I2 =>  inp_feat(135), I3 =>  inp_feat(210), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_0_L_3_inst : LUT6 generic map(INIT => "1000001011111111000011101011100010111010111111111110101111110010") port map( O =>C_43_S_0_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(123), I2 =>  inp_feat(108), I3 =>  inp_feat(248), I4 =>  inp_feat(442), I5 =>  inp_feat(94)); 
C_43_S_0_L_4_inst : LUT6 generic map(INIT => "0000001000111010101000101011100011111111111100000011101011111011") port map( O =>C_43_S_0_L_4_out, I0 =>  inp_feat(182), I1 =>  inp_feat(334), I2 =>  inp_feat(35), I3 =>  inp_feat(282), I4 =>  inp_feat(248), I5 =>  inp_feat(94)); 
C_43_S_0_L_5_inst : LUT6 generic map(INIT => "1101110100101100100111011111111011111111111011001110111000001000") port map( O =>C_43_S_0_L_5_out, I0 =>  inp_feat(300), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_1_L_0_inst : LUT6 generic map(INIT => "1111111010111111111111101110000000100000001111001110100010000000") port map( O =>C_43_S_1_L_0_out, I0 =>  inp_feat(120), I1 =>  inp_feat(381), I2 =>  inp_feat(210), I3 =>  inp_feat(487), I4 =>  inp_feat(434), I5 =>  inp_feat(91)); 
C_43_S_1_L_1_inst : LUT6 generic map(INIT => "0000110111011101111101111101010011111111110111101111110000001100") port map( O =>C_43_S_1_L_1_out, I0 =>  inp_feat(228), I1 =>  inp_feat(470), I2 =>  inp_feat(135), I3 =>  inp_feat(210), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_1_L_2_inst : LUT6 generic map(INIT => "1000001011111111000011101011100010111010111111111110101111110010") port map( O =>C_43_S_1_L_2_out, I0 =>  inp_feat(1), I1 =>  inp_feat(123), I2 =>  inp_feat(108), I3 =>  inp_feat(248), I4 =>  inp_feat(442), I5 =>  inp_feat(94)); 
C_43_S_1_L_3_inst : LUT6 generic map(INIT => "0000001000111010101000101011100011111111111100000011101011111011") port map( O =>C_43_S_1_L_3_out, I0 =>  inp_feat(182), I1 =>  inp_feat(334), I2 =>  inp_feat(35), I3 =>  inp_feat(282), I4 =>  inp_feat(248), I5 =>  inp_feat(94)); 
C_43_S_1_L_4_inst : LUT6 generic map(INIT => "1101110100101100100111011111111011111111111011001110111000001000") port map( O =>C_43_S_1_L_4_out, I0 =>  inp_feat(300), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_1_L_5_inst : LUT6 generic map(INIT => "0010101010011110111111101110101011111111110111001110101000001000") port map( O =>C_43_S_1_L_5_out, I0 =>  inp_feat(209), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_2_L_0_inst : LUT6 generic map(INIT => "1001010100101100100111011111111011111111111011001110111000001000") port map( O =>C_43_S_2_L_0_out, I0 =>  inp_feat(300), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_2_L_1_inst : LUT6 generic map(INIT => "1010101010001101101111001001101011111111111011101111101000000000") port map( O =>C_43_S_2_L_1_out, I0 =>  inp_feat(182), I1 =>  inp_feat(263), I2 =>  inp_feat(61), I3 =>  inp_feat(210), I4 =>  inp_feat(487), I5 =>  inp_feat(434)); 
C_43_S_2_L_2_inst : LUT6 generic map(INIT => "0010010101010101101011011100111111111111111011101111101000000000") port map( O =>C_43_S_2_L_2_out, I0 =>  inp_feat(174), I1 =>  inp_feat(263), I2 =>  inp_feat(61), I3 =>  inp_feat(210), I4 =>  inp_feat(487), I5 =>  inp_feat(434)); 
C_43_S_2_L_3_inst : LUT6 generic map(INIT => "0011100001011111000100000011000111111011111101110111000011110101") port map( O =>C_43_S_2_L_3_out, I0 =>  inp_feat(282), I1 =>  inp_feat(476), I2 =>  inp_feat(25), I3 =>  inp_feat(266), I4 =>  inp_feat(1), I5 =>  inp_feat(94)); 
C_43_S_2_L_4_inst : LUT6 generic map(INIT => "1011001111101110111110100111110011111110111010101011101000100000") port map( O =>C_43_S_2_L_4_out, I0 =>  inp_feat(306), I1 =>  inp_feat(248), I2 =>  inp_feat(184), I3 =>  inp_feat(210), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_2_L_5_inst : LUT6 generic map(INIT => "0010100100011100101111101010111011111111111011001110111000001000") port map( O =>C_43_S_2_L_5_out, I0 =>  inp_feat(213), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_3_L_0_inst : LUT6 generic map(INIT => "1110101000101101011011101101111011111111101011001111111000001000") port map( O =>C_43_S_3_L_0_out, I0 =>  inp_feat(361), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_3_L_1_inst : LUT6 generic map(INIT => "0011100100101010111111101111101111111111111010001100010000000000") port map( O =>C_43_S_3_L_1_out, I0 =>  inp_feat(263), I1 =>  inp_feat(481), I2 =>  inp_feat(429), I3 =>  inp_feat(210), I4 =>  inp_feat(487), I5 =>  inp_feat(434)); 
C_43_S_3_L_2_inst : LUT6 generic map(INIT => "1100110111011110111111010100110011111111111011001110110010110000") port map( O =>C_43_S_3_L_2_out, I0 =>  inp_feat(228), I1 =>  inp_feat(120), I2 =>  inp_feat(42), I3 =>  inp_feat(210), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_3_L_3_inst : LUT6 generic map(INIT => "1000100111011100111111011101110011101100100010001100100000001000") port map( O =>C_43_S_3_L_3_out, I0 =>  inp_feat(106), I1 =>  inp_feat(21), I2 =>  inp_feat(135), I3 =>  inp_feat(210), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_3_L_4_inst : LUT6 generic map(INIT => "1110100010010010111001111010000000001000100000000011100011101000") port map( O =>C_43_S_3_L_4_out, I0 =>  inp_feat(21), I1 =>  inp_feat(488), I2 =>  inp_feat(384), I3 =>  inp_feat(230), I4 =>  inp_feat(395), I5 =>  inp_feat(182)); 
C_43_S_3_L_5_inst : LUT6 generic map(INIT => "0001111101011111000111000101110111111111111111100011110111111111") port map( O =>C_43_S_3_L_5_out, I0 =>  inp_feat(108), I1 =>  inp_feat(479), I2 =>  inp_feat(163), I3 =>  inp_feat(356), I4 =>  inp_feat(114), I5 =>  inp_feat(187)); 
C_43_S_4_L_0_inst : LUT6 generic map(INIT => "1011100110111011011000111111111111111111111010101110111010000000") port map( O =>C_43_S_4_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(228), I2 =>  inp_feat(25), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_4_L_1_inst : LUT6 generic map(INIT => "1011001010110010111010101100111011111111111010111010101010100000") port map( O =>C_43_S_4_L_1_out, I0 =>  inp_feat(399), I1 =>  inp_feat(334), I2 =>  inp_feat(25), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_4_L_2_inst : LUT6 generic map(INIT => "1100110111000100111111101110000111011001000001000010110001110101") port map( O =>C_43_S_4_L_2_out, I0 =>  inp_feat(176), I1 =>  inp_feat(292), I2 =>  inp_feat(494), I3 =>  inp_feat(142), I4 =>  inp_feat(209), I5 =>  inp_feat(232)); 
C_43_S_4_L_3_inst : LUT6 generic map(INIT => "0001010100001000100111011110111111111111111111111110111100000000") port map( O =>C_43_S_4_L_3_out, I0 =>  inp_feat(509), I1 =>  inp_feat(263), I2 =>  inp_feat(61), I3 =>  inp_feat(210), I4 =>  inp_feat(487), I5 =>  inp_feat(434)); 
C_43_S_4_L_4_inst : LUT6 generic map(INIT => "1100011001011001011001101101111111111111110011101100101000000000") port map( O =>C_43_S_4_L_4_out, I0 =>  inp_feat(178), I1 =>  inp_feat(429), I2 =>  inp_feat(61), I3 =>  inp_feat(210), I4 =>  inp_feat(487), I5 =>  inp_feat(434)); 
C_43_S_4_L_5_inst : LUT6 generic map(INIT => "1101011011111010010111001110010011111110111011101111111011100100") port map( O =>C_43_S_4_L_5_out, I0 =>  inp_feat(371), I1 =>  inp_feat(507), I2 =>  inp_feat(234), I3 =>  inp_feat(98), I4 =>  inp_feat(207), I5 =>  inp_feat(51)); 
C_43_S_5_L_0_inst : LUT6 generic map(INIT => "0010111000011110001111101110101011111111110111001110101000001000") port map( O =>C_43_S_5_L_0_out, I0 =>  inp_feat(209), I1 =>  inp_feat(285), I2 =>  inp_feat(490), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_5_L_1_inst : LUT6 generic map(INIT => "0111110101011101011111101000100011111111111111111110101010000000") port map( O =>C_43_S_5_L_1_out, I0 =>  inp_feat(92), I1 =>  inp_feat(418), I2 =>  inp_feat(323), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_5_L_2_inst : LUT6 generic map(INIT => "1110111111110101110010001101100011111111110111011111110111010100") port map( O =>C_43_S_5_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(507), I2 =>  inp_feat(234), I3 =>  inp_feat(98), I4 =>  inp_feat(207), I5 =>  inp_feat(51)); 
C_43_S_5_L_3_inst : LUT6 generic map(INIT => "0001011011101000010011001110010011111111111111101110111011100100") port map( O =>C_43_S_5_L_3_out, I0 =>  inp_feat(371), I1 =>  inp_feat(494), I2 =>  inp_feat(234), I3 =>  inp_feat(98), I4 =>  inp_feat(207), I5 =>  inp_feat(51)); 
C_43_S_5_L_4_inst : LUT6 generic map(INIT => "1110101110011111011110111010001011111111111110111111111100100000") port map( O =>C_43_S_5_L_4_out, I0 =>  inp_feat(62), I1 =>  inp_feat(374), I2 =>  inp_feat(100), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_43_S_5_L_5_inst : LUT6 generic map(INIT => "0011110001111110111011111000100011101111101010001110110010000000") port map( O =>C_43_S_5_L_5_out, I0 =>  inp_feat(10), I1 =>  inp_feat(92), I2 =>  inp_feat(100), I3 =>  inp_feat(487), I4 =>  inp_feat(416), I5 =>  inp_feat(434)); 
C_44_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000") port map( O =>C_44_S_0_L_0_out, I0 =>  inp_feat(453), I1 =>  inp_feat(234), I2 =>  inp_feat(306), I3 =>  inp_feat(10), I4 =>  inp_feat(182), I5 =>  inp_feat(285)); 
C_44_S_0_L_1_inst : LUT6 generic map(INIT => "1110111110101011001010100010111000001000010111100000001000001111") port map( O =>C_44_S_0_L_1_out, I0 =>  inp_feat(403), I1 =>  inp_feat(151), I2 =>  inp_feat(492), I3 =>  inp_feat(371), I4 =>  inp_feat(489), I5 =>  inp_feat(91)); 
C_44_S_0_L_2_inst : LUT6 generic map(INIT => "1110100011111111100010101111111000011110101010000000000000000000") port map( O =>C_44_S_0_L_2_out, I0 =>  inp_feat(306), I1 =>  inp_feat(380), I2 =>  inp_feat(422), I3 =>  inp_feat(391), I4 =>  inp_feat(182), I5 =>  inp_feat(499)); 
C_44_S_0_L_3_inst : LUT6 generic map(INIT => "0101001011110010111100101010111000000010100000001110101110100010") port map( O =>C_44_S_0_L_3_out, I0 =>  inp_feat(91), I1 =>  inp_feat(379), I2 =>  inp_feat(494), I3 =>  inp_feat(98), I4 =>  inp_feat(418), I5 =>  inp_feat(405)); 
C_44_S_0_L_4_inst : LUT6 generic map(INIT => "1100100000011100111111101111111101000000110001000110100011111101") port map( O =>C_44_S_0_L_4_out, I0 =>  inp_feat(378), I1 =>  inp_feat(420), I2 =>  inp_feat(154), I3 =>  inp_feat(106), I4 =>  inp_feat(339), I5 =>  inp_feat(377)); 
C_44_S_0_L_5_inst : LUT6 generic map(INIT => "0101000111110000110010001111110101010000111111110000000001001100") port map( O =>C_44_S_0_L_5_out, I0 =>  inp_feat(282), I1 =>  inp_feat(422), I2 =>  inp_feat(44), I3 =>  inp_feat(391), I4 =>  inp_feat(127), I5 =>  inp_feat(161)); 
C_44_S_1_L_0_inst : LUT6 generic map(INIT => "1110111110101011001010100010111000001000010111100000001000001111") port map( O =>C_44_S_1_L_0_out, I0 =>  inp_feat(403), I1 =>  inp_feat(151), I2 =>  inp_feat(492), I3 =>  inp_feat(371), I4 =>  inp_feat(489), I5 =>  inp_feat(91)); 
C_44_S_1_L_1_inst : LUT6 generic map(INIT => "1110100011111111100010101111111000011110101010000000000000000000") port map( O =>C_44_S_1_L_1_out, I0 =>  inp_feat(306), I1 =>  inp_feat(380), I2 =>  inp_feat(422), I3 =>  inp_feat(391), I4 =>  inp_feat(182), I5 =>  inp_feat(499)); 
C_44_S_1_L_2_inst : LUT6 generic map(INIT => "0101001011110010111100101010111000000010100000001110101110100010") port map( O =>C_44_S_1_L_2_out, I0 =>  inp_feat(91), I1 =>  inp_feat(379), I2 =>  inp_feat(494), I3 =>  inp_feat(98), I4 =>  inp_feat(418), I5 =>  inp_feat(405)); 
C_44_S_1_L_3_inst : LUT6 generic map(INIT => "1100100000011100111111101111111101000000110001000110100011111101") port map( O =>C_44_S_1_L_3_out, I0 =>  inp_feat(378), I1 =>  inp_feat(420), I2 =>  inp_feat(154), I3 =>  inp_feat(106), I4 =>  inp_feat(339), I5 =>  inp_feat(377)); 
C_44_S_1_L_4_inst : LUT6 generic map(INIT => "0101000111110000110010001111110101010000111111110000000001001100") port map( O =>C_44_S_1_L_4_out, I0 =>  inp_feat(282), I1 =>  inp_feat(422), I2 =>  inp_feat(44), I3 =>  inp_feat(391), I4 =>  inp_feat(127), I5 =>  inp_feat(161)); 
C_44_S_1_L_5_inst : LUT6 generic map(INIT => "1111011111111111101110111111110001010111000000101111111011011110") port map( O =>C_44_S_1_L_5_out, I0 =>  inp_feat(120), I1 =>  inp_feat(446), I2 =>  inp_feat(200), I3 =>  inp_feat(389), I4 =>  inp_feat(16), I5 =>  inp_feat(369)); 
C_44_S_2_L_0_inst : LUT6 generic map(INIT => "1111111000001110111000101000001010001100001011101000000010001100") port map( O =>C_44_S_2_L_0_out, I0 =>  inp_feat(371), I1 =>  inp_feat(123), I2 =>  inp_feat(144), I3 =>  inp_feat(356), I4 =>  inp_feat(312), I5 =>  inp_feat(91)); 
C_44_S_2_L_1_inst : LUT6 generic map(INIT => "1000110100111110000011001110100010101011111001111110111011101100") port map( O =>C_44_S_2_L_1_out, I0 =>  inp_feat(507), I1 =>  inp_feat(399), I2 =>  inp_feat(485), I3 =>  inp_feat(434), I4 =>  inp_feat(51), I5 =>  inp_feat(391)); 
C_44_S_2_L_2_inst : LUT6 generic map(INIT => "1111010111110000111101000101010100000001111110111111001111110000") port map( O =>C_44_S_2_L_2_out, I0 =>  inp_feat(37), I1 =>  inp_feat(226), I2 =>  inp_feat(182), I3 =>  inp_feat(7), I4 =>  inp_feat(440), I5 =>  inp_feat(217)); 
C_44_S_2_L_3_inst : LUT6 generic map(INIT => "0010001000110101001000100001001011101111111111110011000011110000") port map( O =>C_44_S_2_L_3_out, I0 =>  inp_feat(179), I1 =>  inp_feat(253), I2 =>  inp_feat(480), I3 =>  inp_feat(59), I4 =>  inp_feat(207), I5 =>  inp_feat(282)); 
C_44_S_2_L_4_inst : LUT6 generic map(INIT => "1110101110000010111011111010101000001001000000001110100111111100") port map( O =>C_44_S_2_L_4_out, I0 =>  inp_feat(453), I1 =>  inp_feat(367), I2 =>  inp_feat(299), I3 =>  inp_feat(338), I4 =>  inp_feat(320), I5 =>  inp_feat(24)); 
C_44_S_2_L_5_inst : LUT6 generic map(INIT => "1011001001011000111111101000000011111000100100000100100001000000") port map( O =>C_44_S_2_L_5_out, I0 =>  inp_feat(311), I1 =>  inp_feat(182), I2 =>  inp_feat(272), I3 =>  inp_feat(44), I4 =>  inp_feat(389), I5 =>  inp_feat(161)); 
C_44_S_3_L_0_inst : LUT6 generic map(INIT => "0000010110111110100011001110100010001010111001111110111011101100") port map( O =>C_44_S_3_L_0_out, I0 =>  inp_feat(507), I1 =>  inp_feat(399), I2 =>  inp_feat(485), I3 =>  inp_feat(434), I4 =>  inp_feat(51), I5 =>  inp_feat(391)); 
C_44_S_3_L_1_inst : LUT6 generic map(INIT => "1111100111110111111111111111111101100100111101101111111101101111") port map( O =>C_44_S_3_L_1_out, I0 =>  inp_feat(11), I1 =>  inp_feat(251), I2 =>  inp_feat(306), I3 =>  inp_feat(19), I4 =>  inp_feat(327), I5 =>  inp_feat(197)); 
C_44_S_3_L_2_inst : LUT6 generic map(INIT => "1100010000110100111101011011000000001101110010000100101011110010") port map( O =>C_44_S_3_L_2_out, I0 =>  inp_feat(71), I1 =>  inp_feat(399), I2 =>  inp_feat(494), I3 =>  inp_feat(332), I4 =>  inp_feat(339), I5 =>  inp_feat(377)); 
C_44_S_3_L_3_inst : LUT6 generic map(INIT => "1011111100100010001000111110101000111010100010000001111111011000") port map( O =>C_44_S_3_L_3_out, I0 =>  inp_feat(207), I1 =>  inp_feat(42), I2 =>  inp_feat(415), I3 =>  inp_feat(405), I4 =>  inp_feat(350), I5 =>  inp_feat(220)); 
C_44_S_3_L_4_inst : LUT6 generic map(INIT => "0101011100111000101111011111000000011111111000001111101110000000") port map( O =>C_44_S_3_L_4_out, I0 =>  inp_feat(404), I1 =>  inp_feat(197), I2 =>  inp_feat(473), I3 =>  inp_feat(363), I4 =>  inp_feat(258), I5 =>  inp_feat(472)); 
C_44_S_3_L_5_inst : LUT6 generic map(INIT => "1101111101100101111110111111010001110110111100101111111100110000") port map( O =>C_44_S_3_L_5_out, I0 =>  inp_feat(156), I1 =>  inp_feat(25), I2 =>  inp_feat(403), I3 =>  inp_feat(122), I4 =>  inp_feat(446), I5 =>  inp_feat(472)); 
C_44_S_4_L_0_inst : LUT6 generic map(INIT => "1111000011111100101100100011001100001000101100011011010110111011") port map( O =>C_44_S_4_L_0_out, I0 =>  inp_feat(17), I1 =>  inp_feat(373), I2 =>  inp_feat(63), I3 =>  inp_feat(467), I4 =>  inp_feat(106), I5 =>  inp_feat(350)); 
C_44_S_4_L_1_inst : LUT6 generic map(INIT => "0101000001111011011111111001001101001100111110011101010100111011") port map( O =>C_44_S_4_L_1_out, I0 =>  inp_feat(445), I1 =>  inp_feat(318), I2 =>  inp_feat(133), I3 =>  inp_feat(266), I4 =>  inp_feat(339), I5 =>  inp_feat(377)); 
C_44_S_4_L_2_inst : LUT6 generic map(INIT => "1000000110011101101110011001010011111111111011001110110001101000") port map( O =>C_44_S_4_L_2_out, I0 =>  inp_feat(132), I1 =>  inp_feat(182), I2 =>  inp_feat(371), I3 =>  inp_feat(44), I4 =>  inp_feat(75), I5 =>  inp_feat(428)); 
C_44_S_4_L_3_inst : LUT6 generic map(INIT => "1111111110011011111010101110001000101011001100101111011111111111") port map( O =>C_44_S_4_L_3_out, I0 =>  inp_feat(71), I1 =>  inp_feat(383), I2 =>  inp_feat(13), I3 =>  inp_feat(106), I4 =>  inp_feat(481), I5 =>  inp_feat(405)); 
C_44_S_4_L_4_inst : LUT6 generic map(INIT => "1101101001000000111011101111111001100000000000001111111111111010") port map( O =>C_44_S_4_L_4_out, I0 =>  inp_feat(162), I1 =>  inp_feat(446), I2 =>  inp_feat(389), I3 =>  inp_feat(413), I4 =>  inp_feat(16), I5 =>  inp_feat(472)); 
C_44_S_4_L_5_inst : LUT6 generic map(INIT => "0001011101110110001111110101111011101111010011111101101001001111") port map( O =>C_44_S_4_L_5_out, I0 =>  inp_feat(130), I1 =>  inp_feat(252), I2 =>  inp_feat(324), I3 =>  inp_feat(311), I4 =>  inp_feat(483), I5 =>  inp_feat(387)); 
C_44_S_5_L_0_inst : LUT6 generic map(INIT => "1010101111011011111011111010001000011011001000101111111110100000") port map( O =>C_44_S_5_L_0_out, I0 =>  inp_feat(10), I1 =>  inp_feat(395), I2 =>  inp_feat(234), I3 =>  inp_feat(306), I4 =>  inp_feat(38), I5 =>  inp_feat(387)); 
C_44_S_5_L_1_inst : LUT6 generic map(INIT => "1100101001011100111111111111111100100000101010001111110011110010") port map( O =>C_44_S_5_L_1_out, I0 =>  inp_feat(72), I1 =>  inp_feat(436), I2 =>  inp_feat(366), I3 =>  inp_feat(416), I4 =>  inp_feat(339), I5 =>  inp_feat(377)); 
C_44_S_5_L_2_inst : LUT6 generic map(INIT => "0011000111100100001110111000100000110010110011101111000000000000") port map( O =>C_44_S_5_L_2_out, I0 =>  inp_feat(142), I1 =>  inp_feat(404), I2 =>  inp_feat(91), I3 =>  inp_feat(193), I4 =>  inp_feat(23), I5 =>  inp_feat(197)); 
C_44_S_5_L_3_inst : LUT6 generic map(INIT => "0101010111101110110101111110111001011100111111100000010011111100") port map( O =>C_44_S_5_L_3_out, I0 =>  inp_feat(344), I1 =>  inp_feat(392), I2 =>  inp_feat(476), I3 =>  inp_feat(445), I4 =>  inp_feat(23), I5 =>  inp_feat(264)); 
C_44_S_5_L_4_inst : LUT6 generic map(INIT => "1100000011101010000000101110110011111111111111111111111111110111") port map( O =>C_44_S_5_L_4_out, I0 =>  inp_feat(207), I1 =>  inp_feat(231), I2 =>  inp_feat(220), I3 =>  inp_feat(336), I4 =>  inp_feat(172), I5 =>  inp_feat(362)); 
C_44_S_5_L_5_inst : LUT6 generic map(INIT => "1001001010011010111110110011111000110011011011111101000000101000") port map( O =>C_44_S_5_L_5_out, I0 =>  inp_feat(377), I1 =>  inp_feat(25), I2 =>  inp_feat(479), I3 =>  inp_feat(120), I4 =>  inp_feat(193), I5 =>  inp_feat(267)); 
C_45_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000000000011100000001000100110001001101111111") port map( O =>C_45_S_0_L_0_out, I0 =>  inp_feat(91), I1 =>  inp_feat(234), I2 =>  inp_feat(306), I3 =>  inp_feat(10), I4 =>  inp_feat(182), I5 =>  inp_feat(285)); 
C_45_S_0_L_1_inst : LUT6 generic map(INIT => "0001000011010101000000000000001010110111111101110000000000000001") port map( O =>C_45_S_0_L_1_out, I0 =>  inp_feat(10), I1 =>  inp_feat(494), I2 =>  inp_feat(175), I3 =>  inp_feat(399), I4 =>  inp_feat(74), I5 =>  inp_feat(123)); 
C_45_S_0_L_2_inst : LUT6 generic map(INIT => "0000000100000111110100110111111110110111010011111001001101110111") port map( O =>C_45_S_0_L_2_out, I0 =>  inp_feat(494), I1 =>  inp_feat(123), I2 =>  inp_feat(272), I3 =>  inp_feat(285), I4 =>  inp_feat(142), I5 =>  inp_feat(279)); 
C_45_S_0_L_3_inst : LUT6 generic map(INIT => "0000000000010000001000101010001000000001110111101010000010111000") port map( O =>C_45_S_0_L_3_out, I0 =>  inp_feat(226), I1 =>  inp_feat(284), I2 =>  inp_feat(395), I3 =>  inp_feat(394), I4 =>  inp_feat(91), I5 =>  inp_feat(359)); 
C_45_S_0_L_4_inst : LUT6 generic map(INIT => "0001100100001100110101110000000011010001100011000101011100000000") port map( O =>C_45_S_0_L_4_out, I0 =>  inp_feat(234), I1 =>  inp_feat(312), I2 =>  inp_feat(182), I3 =>  inp_feat(248), I4 =>  inp_feat(285), I5 =>  inp_feat(461)); 
C_45_S_0_L_5_inst : LUT6 generic map(INIT => "1111000000000001000000010001111100000000000000000000000000010111") port map( O =>C_45_S_0_L_5_out, I0 =>  inp_feat(44), I1 =>  inp_feat(83), I2 =>  inp_feat(226), I3 =>  inp_feat(266), I4 =>  inp_feat(173), I5 =>  inp_feat(293)); 
C_45_S_1_L_0_inst : LUT6 generic map(INIT => "0001000011010101000000000000001010110111111101110000000000000001") port map( O =>C_45_S_1_L_0_out, I0 =>  inp_feat(10), I1 =>  inp_feat(494), I2 =>  inp_feat(175), I3 =>  inp_feat(399), I4 =>  inp_feat(74), I5 =>  inp_feat(123)); 
C_45_S_1_L_1_inst : LUT6 generic map(INIT => "0000000100000111110100110111111110110111010011111001001101110111") port map( O =>C_45_S_1_L_1_out, I0 =>  inp_feat(494), I1 =>  inp_feat(123), I2 =>  inp_feat(272), I3 =>  inp_feat(285), I4 =>  inp_feat(142), I5 =>  inp_feat(279)); 
C_45_S_1_L_2_inst : LUT6 generic map(INIT => "0000000000010000001000101010001000000001110111101010000010111000") port map( O =>C_45_S_1_L_2_out, I0 =>  inp_feat(226), I1 =>  inp_feat(284), I2 =>  inp_feat(395), I3 =>  inp_feat(394), I4 =>  inp_feat(91), I5 =>  inp_feat(359)); 
C_45_S_1_L_3_inst : LUT6 generic map(INIT => "0001100100001100110101110000000011010001100011000101011100000000") port map( O =>C_45_S_1_L_3_out, I0 =>  inp_feat(234), I1 =>  inp_feat(312), I2 =>  inp_feat(182), I3 =>  inp_feat(248), I4 =>  inp_feat(285), I5 =>  inp_feat(461)); 
C_45_S_1_L_4_inst : LUT6 generic map(INIT => "1111000000000001000000010001111100000000000000000000000000010111") port map( O =>C_45_S_1_L_4_out, I0 =>  inp_feat(44), I1 =>  inp_feat(83), I2 =>  inp_feat(226), I3 =>  inp_feat(266), I4 =>  inp_feat(173), I5 =>  inp_feat(293)); 
C_45_S_1_L_5_inst : LUT6 generic map(INIT => "0101010001010101000000000000001011011101111111110000000110000000") port map( O =>C_45_S_1_L_5_out, I0 =>  inp_feat(142), I1 =>  inp_feat(490), I2 =>  inp_feat(292), I3 =>  inp_feat(399), I4 =>  inp_feat(474), I5 =>  inp_feat(454)); 
C_45_S_2_L_0_inst : LUT6 generic map(INIT => "0001000100000000111101110000000110011000000000001111000100000010") port map( O =>C_45_S_2_L_0_out, I0 =>  inp_feat(231), I1 =>  inp_feat(292), I2 =>  inp_feat(472), I3 =>  inp_feat(474), I4 =>  inp_feat(142), I5 =>  inp_feat(226)); 
C_45_S_2_L_1_inst : LUT6 generic map(INIT => "0010110001100010000010010010000011101110011000110010000001100010") port map( O =>C_45_S_2_L_1_out, I0 =>  inp_feat(324), I1 =>  inp_feat(507), I2 =>  inp_feat(168), I3 =>  inp_feat(269), I4 =>  inp_feat(260), I5 =>  inp_feat(231)); 
C_45_S_2_L_2_inst : LUT6 generic map(INIT => "1011011110000101000101010000110100000000000000000000000011000000") port map( O =>C_45_S_2_L_2_out, I0 =>  inp_feat(266), I1 =>  inp_feat(418), I2 =>  inp_feat(476), I3 =>  inp_feat(105), I4 =>  inp_feat(411), I5 =>  inp_feat(183)); 
C_45_S_2_L_3_inst : LUT6 generic map(INIT => "0000000000011110001011010000110000000000001100001100111011101111") port map( O =>C_45_S_2_L_3_out, I0 =>  inp_feat(389), I1 =>  inp_feat(399), I2 =>  inp_feat(418), I3 =>  inp_feat(233), I4 =>  inp_feat(279), I5 =>  inp_feat(180)); 
C_45_S_2_L_4_inst : LUT6 generic map(INIT => "0001000001010010010100001001100011110100011101001101000001011000") port map( O =>C_45_S_2_L_4_out, I0 =>  inp_feat(182), I1 =>  inp_feat(499), I2 =>  inp_feat(368), I3 =>  inp_feat(142), I4 =>  inp_feat(291), I5 =>  inp_feat(196)); 
C_45_S_2_L_5_inst : LUT6 generic map(INIT => "0001010100000010110111110000000010101110000000000000000000000000") port map( O =>C_45_S_2_L_5_out, I0 =>  inp_feat(20), I1 =>  inp_feat(290), I2 =>  inp_feat(429), I3 =>  inp_feat(12), I4 =>  inp_feat(387), I5 =>  inp_feat(263)); 
C_45_S_3_L_0_inst : LUT6 generic map(INIT => "0000010000000011000100001101000110001000101100011101000011110111") port map( O =>C_45_S_3_L_0_out, I0 =>  inp_feat(182), I1 =>  inp_feat(430), I2 =>  inp_feat(133), I3 =>  inp_feat(507), I4 =>  inp_feat(20), I5 =>  inp_feat(231)); 
C_45_S_3_L_1_inst : LUT6 generic map(INIT => "1111010110100010101110011010000000000000000000000000000010000000") port map( O =>C_45_S_3_L_1_out, I0 =>  inp_feat(318), I1 =>  inp_feat(16), I2 =>  inp_feat(441), I3 =>  inp_feat(105), I4 =>  inp_feat(411), I5 =>  inp_feat(183)); 
C_45_S_3_L_2_inst : LUT6 generic map(INIT => "0010001001000101000000000000010000000000000000000000000000000000") port map( O =>C_45_S_3_L_2_out, I0 =>  inp_feat(108), I1 =>  inp_feat(123), I2 =>  inp_feat(282), I3 =>  inp_feat(173), I4 =>  inp_feat(293), I5 =>  inp_feat(14)); 
C_45_S_3_L_3_inst : LUT6 generic map(INIT => "0000110011000000010000000010000011000011000001000111000010010001") port map( O =>C_45_S_3_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(135), I2 =>  inp_feat(316), I3 =>  inp_feat(254), I4 =>  inp_feat(338), I5 =>  inp_feat(415)); 
C_45_S_3_L_4_inst : LUT6 generic map(INIT => "0001100001110011111001000010001000000000000000100110010000100010") port map( O =>C_45_S_3_L_4_out, I0 =>  inp_feat(10), I1 =>  inp_feat(395), I2 =>  inp_feat(105), I3 =>  inp_feat(108), I4 =>  inp_feat(182), I5 =>  inp_feat(3)); 
C_45_S_3_L_5_inst : LUT6 generic map(INIT => "0100101000010000000001000111110010111011110100110000001000000000") port map( O =>C_45_S_3_L_5_out, I0 =>  inp_feat(73), I1 =>  inp_feat(272), I2 =>  inp_feat(142), I3 =>  inp_feat(338), I4 =>  inp_feat(45), I5 =>  inp_feat(479)); 
C_45_S_4_L_0_inst : LUT6 generic map(INIT => "0001001100011101111110110111001110110011000110111111001111110011") port map( O =>C_45_S_4_L_0_out, I0 =>  inp_feat(21), I1 =>  inp_feat(494), I2 =>  inp_feat(478), I3 =>  inp_feat(196), I4 =>  inp_feat(91), I5 =>  inp_feat(126)); 
C_45_S_4_L_1_inst : LUT6 generic map(INIT => "0010101010001010000100101010000001100010100000100000001001010010") port map( O =>C_45_S_4_L_1_out, I0 =>  inp_feat(248), I1 =>  inp_feat(91), I2 =>  inp_feat(498), I3 =>  inp_feat(250), I4 =>  inp_feat(83), I5 =>  inp_feat(461)); 
C_45_S_4_L_2_inst : LUT6 generic map(INIT => "1001001100011010010000001000000000000000010000001000000000000000") port map( O =>C_45_S_4_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(377), I2 =>  inp_feat(132), I3 =>  inp_feat(416), I4 =>  inp_feat(226), I5 =>  inp_feat(256)); 
C_45_S_4_L_3_inst : LUT6 generic map(INIT => "1001000100000011010000000000110000000100000011010100111111101110") port map( O =>C_45_S_4_L_3_out, I0 =>  inp_feat(411), I1 =>  inp_feat(327), I2 =>  inp_feat(157), I3 =>  inp_feat(37), I4 =>  inp_feat(282), I5 =>  inp_feat(266)); 
C_45_S_4_L_4_inst : LUT6 generic map(INIT => "0100000000000000000110010000000000000000010000000111000100000100") port map( O =>C_45_S_4_L_4_out, I0 =>  inp_feat(11), I1 =>  inp_feat(321), I2 =>  inp_feat(441), I3 =>  inp_feat(19), I4 =>  inp_feat(417), I5 =>  inp_feat(348)); 
C_45_S_4_L_5_inst : LUT6 generic map(INIT => "0010100100011100100011000100110010010001000000000010101011000010") port map( O =>C_45_S_4_L_5_out, I0 =>  inp_feat(99), I1 =>  inp_feat(510), I2 =>  inp_feat(320), I3 =>  inp_feat(77), I4 =>  inp_feat(157), I5 =>  inp_feat(196)); 
C_45_S_5_L_0_inst : LUT6 generic map(INIT => "0011000111010000111001000000000000000000000000000000000000000000") port map( O =>C_45_S_5_L_0_out, I0 =>  inp_feat(180), I1 =>  inp_feat(184), I2 =>  inp_feat(183), I3 =>  inp_feat(418), I4 =>  inp_feat(292), I5 =>  inp_feat(14)); 
C_45_S_5_L_1_inst : LUT6 generic map(INIT => "1100110010110111000001101011111001000100000100000100010000100100") port map( O =>C_45_S_5_L_1_out, I0 =>  inp_feat(494), I1 =>  inp_feat(248), I2 =>  inp_feat(345), I3 =>  inp_feat(445), I4 =>  inp_feat(151), I5 =>  inp_feat(38)); 
C_45_S_5_L_2_inst : LUT6 generic map(INIT => "0100011000000000000100010000000010010000000000000000000000000001") port map( O =>C_45_S_5_L_2_out, I0 =>  inp_feat(429), I1 =>  inp_feat(176), I2 =>  inp_feat(40), I3 =>  inp_feat(337), I4 =>  inp_feat(423), I5 =>  inp_feat(3)); 
C_45_S_5_L_3_inst : LUT6 generic map(INIT => "0100000000000011110011110000001011010100101101010100000000000001") port map( O =>C_45_S_5_L_3_out, I0 =>  inp_feat(242), I1 =>  inp_feat(389), I2 =>  inp_feat(141), I3 =>  inp_feat(87), I4 =>  inp_feat(231), I5 =>  inp_feat(403)); 
C_45_S_5_L_4_inst : LUT6 generic map(INIT => "0000101100010000110111110000000000000000110000110101011100000000") port map( O =>C_45_S_5_L_4_out, I0 =>  inp_feat(123), I1 =>  inp_feat(250), I2 =>  inp_feat(485), I3 =>  inp_feat(214), I4 =>  inp_feat(272), I5 =>  inp_feat(489)); 
C_45_S_5_L_5_inst : LUT6 generic map(INIT => "1101110101100000001000001111000000000000000010001101000110100000") port map( O =>C_45_S_5_L_5_out, I0 =>  inp_feat(320), I1 =>  inp_feat(207), I2 =>  inp_feat(64), I3 =>  inp_feat(480), I4 =>  inp_feat(175), I5 =>  inp_feat(238)); 
C_46_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111101110100011111110111010001110100010000000") port map( O =>C_46_S_0_L_0_out, I0 =>  inp_feat(453), I1 =>  inp_feat(234), I2 =>  inp_feat(306), I3 =>  inp_feat(10), I4 =>  inp_feat(182), I5 =>  inp_feat(285)); 
C_46_S_0_L_1_inst : LUT6 generic map(INIT => "1110010011100010111001111110111100100000011000001100001011111110") port map( O =>C_46_S_0_L_1_out, I0 =>  inp_feat(20), I1 =>  inp_feat(234), I2 =>  inp_feat(91), I3 =>  inp_feat(413), I4 =>  inp_feat(183), I5 =>  inp_feat(306)); 
C_46_S_0_L_2_inst : LUT6 generic map(INIT => "0010001001111011001000111011001111100001111111110110010111110010") port map( O =>C_46_S_0_L_2_out, I0 =>  inp_feat(20), I1 =>  inp_feat(221), I2 =>  inp_feat(350), I3 =>  inp_feat(45), I4 =>  inp_feat(72), I5 =>  inp_feat(183)); 
C_46_S_0_L_3_inst : LUT6 generic map(INIT => "1010111110101110000011100110111011111011110100110000110011111100") port map( O =>C_46_S_0_L_3_out, I0 =>  inp_feat(350), I1 =>  inp_feat(483), I2 =>  inp_feat(468), I3 =>  inp_feat(222), I4 =>  inp_feat(10), I5 =>  inp_feat(180)); 
C_46_S_0_L_4_inst : LUT6 generic map(INIT => "1001111100101111111111100111111100001100000101101111011001000100") port map( O =>C_46_S_0_L_4_out, I0 =>  inp_feat(283), I1 =>  inp_feat(333), I2 =>  inp_feat(183), I3 =>  inp_feat(32), I4 =>  inp_feat(180), I5 =>  inp_feat(472)); 
C_46_S_0_L_5_inst : LUT6 generic map(INIT => "0101010011111111000111111111101100100001001111100010001100011111") port map( O =>C_46_S_0_L_5_out, I0 =>  inp_feat(483), I1 =>  inp_feat(306), I2 =>  inp_feat(58), I3 =>  inp_feat(416), I4 =>  inp_feat(299), I5 =>  inp_feat(70)); 
C_46_S_1_L_0_inst : LUT6 generic map(INIT => "1110010011100010111001111110111100100000011000001100001011111110") port map( O =>C_46_S_1_L_0_out, I0 =>  inp_feat(20), I1 =>  inp_feat(234), I2 =>  inp_feat(91), I3 =>  inp_feat(413), I4 =>  inp_feat(183), I5 =>  inp_feat(306)); 
C_46_S_1_L_1_inst : LUT6 generic map(INIT => "0010001001111011001000111011001111100001111111110110010111110010") port map( O =>C_46_S_1_L_1_out, I0 =>  inp_feat(20), I1 =>  inp_feat(221), I2 =>  inp_feat(350), I3 =>  inp_feat(45), I4 =>  inp_feat(72), I5 =>  inp_feat(183)); 
C_46_S_1_L_2_inst : LUT6 generic map(INIT => "1010111110101110000011100110111011111011110100110000110011111100") port map( O =>C_46_S_1_L_2_out, I0 =>  inp_feat(350), I1 =>  inp_feat(483), I2 =>  inp_feat(468), I3 =>  inp_feat(222), I4 =>  inp_feat(10), I5 =>  inp_feat(180)); 
C_46_S_1_L_3_inst : LUT6 generic map(INIT => "1001111100101111111111100111111100001100000101101111011001000100") port map( O =>C_46_S_1_L_3_out, I0 =>  inp_feat(283), I1 =>  inp_feat(333), I2 =>  inp_feat(183), I3 =>  inp_feat(32), I4 =>  inp_feat(180), I5 =>  inp_feat(472)); 
C_46_S_1_L_4_inst : LUT6 generic map(INIT => "0101010011111111000111111111101100100001001111100010001100011111") port map( O =>C_46_S_1_L_4_out, I0 =>  inp_feat(483), I1 =>  inp_feat(306), I2 =>  inp_feat(58), I3 =>  inp_feat(416), I4 =>  inp_feat(299), I5 =>  inp_feat(70)); 
C_46_S_1_L_5_inst : LUT6 generic map(INIT => "1111000111110001010000001010000111111111111111111101111111000110") port map( O =>C_46_S_1_L_5_out, I0 =>  inp_feat(334), I1 =>  inp_feat(355), I2 =>  inp_feat(348), I3 =>  inp_feat(409), I4 =>  inp_feat(203), I5 =>  inp_feat(435)); 
C_46_S_2_L_0_inst : LUT6 generic map(INIT => "0000001011111011000000100011101111111111100111110011111111110011") port map( O =>C_46_S_2_L_0_out, I0 =>  inp_feat(11), I1 =>  inp_feat(334), I2 =>  inp_feat(104), I3 =>  inp_feat(180), I4 =>  inp_feat(399), I5 =>  inp_feat(183)); 
C_46_S_2_L_1_inst : LUT6 generic map(INIT => "1111101011100101001011001100111101001000110100010000000010100000") port map( O =>C_46_S_2_L_1_out, I0 =>  inp_feat(91), I1 =>  inp_feat(231), I2 =>  inp_feat(251), I3 =>  inp_feat(187), I4 =>  inp_feat(311), I5 =>  inp_feat(10)); 
C_46_S_2_L_2_inst : LUT6 generic map(INIT => "0010011111100110000001111110111110011111111110110000011111111111") port map( O =>C_46_S_2_L_2_out, I0 =>  inp_feat(452), I1 =>  inp_feat(181), I2 =>  inp_feat(49), I3 =>  inp_feat(73), I4 =>  inp_feat(315), I5 =>  inp_feat(434)); 
C_46_S_2_L_3_inst : LUT6 generic map(INIT => "1111001100001110101011111000001011011011111110001111111110000000") port map( O =>C_46_S_2_L_3_out, I0 =>  inp_feat(234), I1 =>  inp_feat(285), I2 =>  inp_feat(233), I3 =>  inp_feat(272), I4 =>  inp_feat(44), I5 =>  inp_feat(173)); 
C_46_S_2_L_4_inst : LUT6 generic map(INIT => "1000000010100000010011010110100011111111110010000101111011101000") port map( O =>C_46_S_2_L_4_out, I0 =>  inp_feat(189), I1 =>  inp_feat(217), I2 =>  inp_feat(285), I3 =>  inp_feat(483), I4 =>  inp_feat(456), I5 =>  inp_feat(431)); 
C_46_S_2_L_5_inst : LUT6 generic map(INIT => "0001100011001100000111001001111111101111111111110011010111011111") port map( O =>C_46_S_2_L_5_out, I0 =>  inp_feat(456), I1 =>  inp_feat(70), I2 =>  inp_feat(48), I3 =>  inp_feat(151), I4 =>  inp_feat(348), I5 =>  inp_feat(431)); 
C_46_S_3_L_0_inst : LUT6 generic map(INIT => "0010000111100011001000111111101111111111111101110011001111111010") port map( O =>C_46_S_3_L_0_out, I0 =>  inp_feat(257), I1 =>  inp_feat(87), I2 =>  inp_feat(70), I3 =>  inp_feat(322), I4 =>  inp_feat(315), I5 =>  inp_feat(434)); 
C_46_S_3_L_1_inst : LUT6 generic map(INIT => "1111111010111010001011010111110111111011001011110000000011001000") port map( O =>C_46_S_3_L_1_out, I0 =>  inp_feat(450), I1 =>  inp_feat(332), I2 =>  inp_feat(391), I3 =>  inp_feat(48), I4 =>  inp_feat(371), I5 =>  inp_feat(430)); 
C_46_S_3_L_2_inst : LUT6 generic map(INIT => "1110101011011111101010101101110100011110111111001110000011100000") port map( O =>C_46_S_3_L_2_out, I0 =>  inp_feat(234), I1 =>  inp_feat(480), I2 =>  inp_feat(10), I3 =>  inp_feat(440), I4 =>  inp_feat(499), I5 =>  inp_feat(182)); 
C_46_S_3_L_3_inst : LUT6 generic map(INIT => "0000001100111011010101011101111101010111011111111111111111110011") port map( O =>C_46_S_3_L_3_out, I0 =>  inp_feat(189), I1 =>  inp_feat(42), I2 =>  inp_feat(229), I3 =>  inp_feat(437), I4 =>  inp_feat(395), I5 =>  inp_feat(238)); 
C_46_S_3_L_4_inst : LUT6 generic map(INIT => "0110111111100000111011101000000011101110101011001100111011000100") port map( O =>C_46_S_3_L_4_out, I0 =>  inp_feat(507), I1 =>  inp_feat(488), I2 =>  inp_feat(44), I3 =>  inp_feat(20), I4 =>  inp_feat(259), I5 =>  inp_feat(435)); 
C_46_S_3_L_5_inst : LUT6 generic map(INIT => "1011100110101111110011001100111100000000101101011000110111101111") port map( O =>C_46_S_3_L_5_out, I0 =>  inp_feat(225), I1 =>  inp_feat(378), I2 =>  inp_feat(272), I3 =>  inp_feat(221), I4 =>  inp_feat(204), I5 =>  inp_feat(479)); 
C_46_S_4_L_0_inst : LUT6 generic map(INIT => "0000010111101101111111110011111010101000110111111111111111110000") port map( O =>C_46_S_4_L_0_out, I0 =>  inp_feat(173), I1 =>  inp_feat(75), I2 =>  inp_feat(465), I3 =>  inp_feat(132), I4 =>  inp_feat(151), I5 =>  inp_feat(63)); 
C_46_S_4_L_1_inst : LUT6 generic map(INIT => "0000010111110110000000001110111011111100100111000111000011111000") port map( O =>C_46_S_4_L_1_out, I0 =>  inp_feat(128), I1 =>  inp_feat(442), I2 =>  inp_feat(166), I3 =>  inp_feat(432), I4 =>  inp_feat(347), I5 =>  inp_feat(222)); 
C_46_S_4_L_2_inst : LUT6 generic map(INIT => "1011101001111110010101011111110111110110110111100011001011111110") port map( O =>C_46_S_4_L_2_out, I0 =>  inp_feat(453), I1 =>  inp_feat(485), I2 =>  inp_feat(152), I3 =>  inp_feat(74), I4 =>  inp_feat(373), I5 =>  inp_feat(173)); 
C_46_S_4_L_3_inst : LUT6 generic map(INIT => "0000101010111111100111101111111111111110010111110000110001111111") port map( O =>C_46_S_4_L_3_out, I0 =>  inp_feat(254), I1 =>  inp_feat(32), I2 =>  inp_feat(54), I3 =>  inp_feat(151), I4 =>  inp_feat(208), I5 =>  inp_feat(322)); 
C_46_S_4_L_4_inst : LUT6 generic map(INIT => "1010101101110011101111001111110011101111001010011111111111011011") port map( O =>C_46_S_4_L_4_out, I0 =>  inp_feat(44), I1 =>  inp_feat(114), I2 =>  inp_feat(450), I3 =>  inp_feat(72), I4 =>  inp_feat(202), I5 =>  inp_feat(187)); 
C_46_S_4_L_5_inst : LUT6 generic map(INIT => "0101001110101101111111011111110111011111100001011111111111010111") port map( O =>C_46_S_4_L_5_out, I0 =>  inp_feat(323), I1 =>  inp_feat(114), I2 =>  inp_feat(450), I3 =>  inp_feat(72), I4 =>  inp_feat(202), I5 =>  inp_feat(187)); 
C_46_S_5_L_0_inst : LUT6 generic map(INIT => "0110111101110101111011001111111100000101010101010111111111111101") port map( O =>C_46_S_5_L_0_out, I0 =>  inp_feat(238), I1 =>  inp_feat(278), I2 =>  inp_feat(106), I3 =>  inp_feat(510), I4 =>  inp_feat(108), I5 =>  inp_feat(31)); 
C_46_S_5_L_1_inst : LUT6 generic map(INIT => "0101101100100011011000100111001011111111111111010100110001011101") port map( O =>C_46_S_5_L_1_out, I0 =>  inp_feat(173), I1 =>  inp_feat(221), I2 =>  inp_feat(54), I3 =>  inp_feat(257), I4 =>  inp_feat(218), I5 =>  inp_feat(435)); 
C_46_S_5_L_2_inst : LUT6 generic map(INIT => "1111110111010101100111111101101101011000100000000000000010000000") port map( O =>C_46_S_5_L_2_out, I0 =>  inp_feat(307), I1 =>  inp_feat(182), I2 =>  inp_feat(20), I3 =>  inp_feat(272), I4 =>  inp_feat(373), I5 =>  inp_feat(472)); 
C_46_S_5_L_3_inst : LUT6 generic map(INIT => "0111110011101010011001101100000000011000000011001111100011001000") port map( O =>C_46_S_5_L_3_out, I0 =>  inp_feat(39), I1 =>  inp_feat(231), I2 =>  inp_feat(371), I3 =>  inp_feat(2), I4 =>  inp_feat(87), I5 =>  inp_feat(264)); 
C_46_S_5_L_4_inst : LUT6 generic map(INIT => "1000100111010000010001011011101010101110111111010110001001101110") port map( O =>C_46_S_5_L_4_out, I0 =>  inp_feat(195), I1 =>  inp_feat(466), I2 =>  inp_feat(269), I3 =>  inp_feat(322), I4 =>  inp_feat(13), I5 =>  inp_feat(200)); 
C_46_S_5_L_5_inst : LUT6 generic map(INIT => "0011111101010001011101111101110111111111111110111100010111111111") port map( O =>C_46_S_5_L_5_out, I0 =>  inp_feat(202), I1 =>  inp_feat(303), I2 =>  inp_feat(407), I3 =>  inp_feat(115), I4 =>  inp_feat(479), I5 =>  inp_feat(18)); 
C_47_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000000000011100000001000100110001001101111111") port map( O =>C_47_S_0_L_0_out, I0 =>  inp_feat(91), I1 =>  inp_feat(234), I2 =>  inp_feat(306), I3 =>  inp_feat(10), I4 =>  inp_feat(182), I5 =>  inp_feat(285)); 
C_47_S_0_L_1_inst : LUT6 generic map(INIT => "1100010010010000110000000100000100000000000000000000000010010000") port map( O =>C_47_S_0_L_1_out, I0 =>  inp_feat(33), I1 =>  inp_feat(374), I2 =>  inp_feat(317), I3 =>  inp_feat(107), I4 =>  inp_feat(267), I5 =>  inp_feat(183)); 
C_47_S_0_L_2_inst : LUT6 generic map(INIT => "0001000000000000000000100000100011101010110000000000001010000000") port map( O =>C_47_S_0_L_2_out, I0 =>  inp_feat(130), I1 =>  inp_feat(207), I2 =>  inp_feat(1), I3 =>  inp_feat(233), I4 =>  inp_feat(418), I5 =>  inp_feat(123)); 
C_47_S_0_L_3_inst : LUT6 generic map(INIT => "1110011111111110000000001110000000000110000000010000000000000000") port map( O =>C_47_S_0_L_3_out, I0 =>  inp_feat(407), I1 =>  inp_feat(257), I2 =>  inp_feat(181), I3 =>  inp_feat(403), I4 =>  inp_feat(435), I5 =>  inp_feat(289)); 
C_47_S_0_L_4_inst : LUT6 generic map(INIT => "0111110011100100000000000110000000000000000100101010000000000000") port map( O =>C_47_S_0_L_4_out, I0 =>  inp_feat(126), I1 =>  inp_feat(72), I2 =>  inp_feat(317), I3 =>  inp_feat(33), I4 =>  inp_feat(183), I5 =>  inp_feat(319)); 
C_47_S_0_L_5_inst : LUT6 generic map(INIT => "0000101010101110000000000000100010101110111011110000100000001110") port map( O =>C_47_S_0_L_5_out, I0 =>  inp_feat(254), I1 =>  inp_feat(449), I2 =>  inp_feat(269), I3 =>  inp_feat(24), I4 =>  inp_feat(104), I5 =>  inp_feat(483)); 
C_47_S_1_L_0_inst : LUT6 generic map(INIT => "1100010010010000110000000100000100000000000000000000000010010000") port map( O =>C_47_S_1_L_0_out, I0 =>  inp_feat(33), I1 =>  inp_feat(374), I2 =>  inp_feat(317), I3 =>  inp_feat(107), I4 =>  inp_feat(267), I5 =>  inp_feat(183)); 
C_47_S_1_L_1_inst : LUT6 generic map(INIT => "0001000000000000000000100000100011101010110000000000001010000000") port map( O =>C_47_S_1_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(207), I2 =>  inp_feat(1), I3 =>  inp_feat(233), I4 =>  inp_feat(418), I5 =>  inp_feat(123)); 
C_47_S_1_L_2_inst : LUT6 generic map(INIT => "1110011111111110000000001110000000000110000000010000000000000000") port map( O =>C_47_S_1_L_2_out, I0 =>  inp_feat(407), I1 =>  inp_feat(257), I2 =>  inp_feat(181), I3 =>  inp_feat(403), I4 =>  inp_feat(435), I5 =>  inp_feat(289)); 
C_47_S_1_L_3_inst : LUT6 generic map(INIT => "0111110011100100000000000110000000000000000100101010000000000000") port map( O =>C_47_S_1_L_3_out, I0 =>  inp_feat(126), I1 =>  inp_feat(72), I2 =>  inp_feat(317), I3 =>  inp_feat(33), I4 =>  inp_feat(183), I5 =>  inp_feat(319)); 
C_47_S_1_L_4_inst : LUT6 generic map(INIT => "0000101010101110000000000000100010101110111011110000100000001110") port map( O =>C_47_S_1_L_4_out, I0 =>  inp_feat(254), I1 =>  inp_feat(449), I2 =>  inp_feat(269), I3 =>  inp_feat(24), I4 =>  inp_feat(104), I5 =>  inp_feat(483)); 
C_47_S_1_L_5_inst : LUT6 generic map(INIT => "1111010001001100101001010010000001100110000000100000000000001100") port map( O =>C_47_S_1_L_5_out, I0 =>  inp_feat(92), I1 =>  inp_feat(464), I2 =>  inp_feat(33), I3 =>  inp_feat(46), I4 =>  inp_feat(288), I5 =>  inp_feat(484)); 
C_47_S_2_L_0_inst : LUT6 generic map(INIT => "0000111110111010111000000100001000000001000000000000010010000000") port map( O =>C_47_S_2_L_0_out, I0 =>  inp_feat(33), I1 =>  inp_feat(244), I2 =>  inp_feat(510), I3 =>  inp_feat(224), I4 =>  inp_feat(267), I5 =>  inp_feat(183)); 
C_47_S_2_L_1_inst : LUT6 generic map(INIT => "0101010100000010000001100010000000000011000000000000001000000000") port map( O =>C_47_S_2_L_1_out, I0 =>  inp_feat(24), I1 =>  inp_feat(140), I2 =>  inp_feat(33), I3 =>  inp_feat(183), I4 =>  inp_feat(319), I5 =>  inp_feat(484)); 
C_47_S_2_L_2_inst : LUT6 generic map(INIT => "1011101000110000100110000000100000111100000001000000000001010000") port map( O =>C_47_S_2_L_2_out, I0 =>  inp_feat(33), I1 =>  inp_feat(92), I2 =>  inp_feat(464), I3 =>  inp_feat(46), I4 =>  inp_feat(288), I5 =>  inp_feat(484)); 
C_47_S_2_L_3_inst : LUT6 generic map(INIT => "0111011000001000011100010000000000010001000000000000000000001000") port map( O =>C_47_S_2_L_3_out, I0 =>  inp_feat(44), I1 =>  inp_feat(94), I2 =>  inp_feat(95), I3 =>  inp_feat(45), I4 =>  inp_feat(435), I5 =>  inp_feat(418)); 
C_47_S_2_L_4_inst : LUT6 generic map(INIT => "0001101001110000000100100000000011111101111100100001000001100000") port map( O =>C_47_S_2_L_4_out, I0 =>  inp_feat(420), I1 =>  inp_feat(181), I2 =>  inp_feat(453), I3 =>  inp_feat(263), I4 =>  inp_feat(289), I5 =>  inp_feat(136)); 
C_47_S_2_L_5_inst : LUT6 generic map(INIT => "1011101110011000111110000000100000000011000000000000000000010001") port map( O =>C_47_S_2_L_5_out, I0 =>  inp_feat(261), I1 =>  inp_feat(456), I2 =>  inp_feat(182), I3 =>  inp_feat(375), I4 =>  inp_feat(6), I5 =>  inp_feat(434)); 
C_47_S_3_L_0_inst : LUT6 generic map(INIT => "0001100100011000111110000000100000000011000000000000000000010001") port map( O =>C_47_S_3_L_0_out, I0 =>  inp_feat(261), I1 =>  inp_feat(456), I2 =>  inp_feat(182), I3 =>  inp_feat(375), I4 =>  inp_feat(6), I5 =>  inp_feat(434)); 
C_47_S_3_L_1_inst : LUT6 generic map(INIT => "1110000000010011110110010000001100000000000000000000010000000110") port map( O =>C_47_S_3_L_1_out, I0 =>  inp_feat(329), I1 =>  inp_feat(150), I2 =>  inp_feat(261), I3 =>  inp_feat(491), I4 =>  inp_feat(456), I5 =>  inp_feat(434)); 
C_47_S_3_L_2_inst : LUT6 generic map(INIT => "0001010000000001000101100000000011101110000101101010011100000000") port map( O =>C_47_S_3_L_2_out, I0 =>  inp_feat(59), I1 =>  inp_feat(33), I2 =>  inp_feat(283), I3 =>  inp_feat(296), I4 =>  inp_feat(277), I5 =>  inp_feat(179)); 
C_47_S_3_L_3_inst : LUT6 generic map(INIT => "1110001101000011011011101011011101010101000000000111111000000010") port map( O =>C_47_S_3_L_3_out, I0 =>  inp_feat(207), I1 =>  inp_feat(300), I2 =>  inp_feat(24), I3 =>  inp_feat(449), I4 =>  inp_feat(269), I5 =>  inp_feat(104)); 
C_47_S_3_L_4_inst : LUT6 generic map(INIT => "1101100010000000111100010000000000000100000100001111101100000000") port map( O =>C_47_S_3_L_4_out, I0 =>  inp_feat(70), I1 =>  inp_feat(285), I2 =>  inp_feat(435), I3 =>  inp_feat(418), I4 =>  inp_feat(272), I5 =>  inp_feat(413)); 
C_47_S_3_L_5_inst : LUT6 generic map(INIT => "0001000100000000110010011010010001000010000000011111011100010001") port map( O =>C_47_S_3_L_5_out, I0 =>  inp_feat(465), I1 =>  inp_feat(230), I2 =>  inp_feat(173), I3 =>  inp_feat(218), I4 =>  inp_feat(471), I5 =>  inp_feat(293)); 
C_47_S_4_L_0_inst : LUT6 generic map(INIT => "1101110111010111001000000000000011111011000101110000000000000000") port map( O =>C_47_S_4_L_0_out, I0 =>  inp_feat(272), I1 =>  inp_feat(494), I2 =>  inp_feat(182), I3 =>  inp_feat(61), I4 =>  inp_feat(352), I5 =>  inp_feat(370)); 
C_47_S_4_L_1_inst : LUT6 generic map(INIT => "1101110110110000001110010000100001110001000000010000000000010000") port map( O =>C_47_S_4_L_1_out, I0 =>  inp_feat(140), I1 =>  inp_feat(33), I2 =>  inp_feat(464), I3 =>  inp_feat(46), I4 =>  inp_feat(288), I5 =>  inp_feat(484)); 
C_47_S_4_L_2_inst : LUT6 generic map(INIT => "1000011001011000011000100000100000000000000000000010000000001100") port map( O =>C_47_S_4_L_2_out, I0 =>  inp_feat(362), I1 =>  inp_feat(465), I2 =>  inp_feat(261), I3 =>  inp_feat(491), I4 =>  inp_feat(456), I5 =>  inp_feat(434)); 
C_47_S_4_L_3_inst : LUT6 generic map(INIT => "0000001000010001101000010001000100000000000000000010000000001100") port map( O =>C_47_S_4_L_3_out, I0 =>  inp_feat(482), I1 =>  inp_feat(445), I2 =>  inp_feat(447), I3 =>  inp_feat(491), I4 =>  inp_feat(456), I5 =>  inp_feat(434)); 
C_47_S_4_L_4_inst : LUT6 generic map(INIT => "1010100010100010001000001000000000000000000000000000001100000110") port map( O =>C_47_S_4_L_4_out, I0 =>  inp_feat(476), I1 =>  inp_feat(182), I2 =>  inp_feat(348), I3 =>  inp_feat(6), I4 =>  inp_feat(456), I5 =>  inp_feat(434)); 
C_47_S_4_L_5_inst : LUT6 generic map(INIT => "0001000100010111000100000000000011111001101000010000000000000000") port map( O =>C_47_S_4_L_5_out, I0 =>  inp_feat(123), I1 =>  inp_feat(371), I2 =>  inp_feat(507), I3 =>  inp_feat(301), I4 =>  inp_feat(60), I5 =>  inp_feat(357)); 
C_47_S_5_L_0_inst : LUT6 generic map(INIT => "1111000011010001101100010100001100000000000000000010000000001100") port map( O =>C_47_S_5_L_0_out, I0 =>  inp_feat(380), I1 =>  inp_feat(440), I2 =>  inp_feat(447), I3 =>  inp_feat(491), I4 =>  inp_feat(456), I5 =>  inp_feat(434)); 
C_47_S_5_L_1_inst : LUT6 generic map(INIT => "0010010011001110000001011011101000000000001010000000100111000011") port map( O =>C_47_S_5_L_1_out, I0 =>  inp_feat(212), I1 =>  inp_feat(456), I2 =>  inp_feat(306), I3 =>  inp_feat(237), I4 =>  inp_feat(160), I5 =>  inp_feat(202)); 
C_47_S_5_L_2_inst : LUT6 generic map(INIT => "1001111000101100101001101111100100000000000010000000110011001000") port map( O =>C_47_S_5_L_2_out, I0 =>  inp_feat(145), I1 =>  inp_feat(254), I2 =>  inp_feat(306), I3 =>  inp_feat(237), I4 =>  inp_feat(160), I5 =>  inp_feat(202)); 
C_47_S_5_L_3_inst : LUT6 generic map(INIT => "0000101010001000011000001000000000000000000000101101010010111001") port map( O =>C_47_S_5_L_3_out, I0 =>  inp_feat(223), I1 =>  inp_feat(319), I2 =>  inp_feat(0), I3 =>  inp_feat(336), I4 =>  inp_feat(510), I5 =>  inp_feat(286)); 
C_47_S_5_L_4_inst : LUT6 generic map(INIT => "1101001010011001000000111111011110011001000001010010011101111111") port map( O =>C_47_S_5_L_4_out, I0 =>  inp_feat(454), I1 =>  inp_feat(234), I2 =>  inp_feat(494), I3 =>  inp_feat(507), I4 =>  inp_feat(371), I5 =>  inp_feat(311)); 
C_47_S_5_L_5_inst : LUT6 generic map(INIT => "0000011000100101001101111101011101010101000001010011011100111111") port map( O =>C_47_S_5_L_5_out, I0 =>  inp_feat(91), I1 =>  inp_feat(123), I2 =>  inp_feat(494), I3 =>  inp_feat(20), I4 =>  inp_feat(371), I5 =>  inp_feat(311)); 
C_48_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000010001000000010011011100000000000100010100010101111111") port map( O =>C_48_S_0_L_0_out, I0 =>  inp_feat(246), I1 =>  inp_feat(183), I2 =>  inp_feat(51), I3 =>  inp_feat(378), I4 =>  inp_feat(317), I5 =>  inp_feat(469)); 
C_48_S_0_L_1_inst : LUT6 generic map(INIT => "0001000001110000011000001111001000110001111100011111001011110011") port map( O =>C_48_S_0_L_1_out, I0 =>  inp_feat(74), I1 =>  inp_feat(469), I2 =>  inp_feat(488), I3 =>  inp_feat(208), I4 =>  inp_feat(328), I5 =>  inp_feat(289)); 
C_48_S_0_L_2_inst : LUT6 generic map(INIT => "0001111100000011111111010000011100000000000000000000000010000000") port map( O =>C_48_S_0_L_2_out, I0 =>  inp_feat(51), I1 =>  inp_feat(81), I2 =>  inp_feat(13), I3 =>  inp_feat(167), I4 =>  inp_feat(33), I5 =>  inp_feat(59)); 
C_48_S_0_L_3_inst : LUT6 generic map(INIT => "0000010101000000000000000000000011001101010011000000000000000100") port map( O =>C_48_S_0_L_3_out, I0 =>  inp_feat(249), I1 =>  inp_feat(436), I2 =>  inp_feat(139), I3 =>  inp_feat(15), I4 =>  inp_feat(186), I5 =>  inp_feat(151)); 
C_48_S_0_L_4_inst : LUT6 generic map(INIT => "0110011001100010010100100101001000000000000000000000000000000010") port map( O =>C_48_S_0_L_4_out, I0 =>  inp_feat(33), I1 =>  inp_feat(375), I2 =>  inp_feat(288), I3 =>  inp_feat(192), I4 =>  inp_feat(368), I5 =>  inp_feat(128)); 
C_48_S_0_L_5_inst : LUT6 generic map(INIT => "0100101101100111000100010101110110111111011111110000000101010111") port map( O =>C_48_S_0_L_5_out, I0 =>  inp_feat(246), I1 =>  inp_feat(139), I2 =>  inp_feat(482), I3 =>  inp_feat(149), I4 =>  inp_feat(494), I5 =>  inp_feat(4)); 
C_48_S_1_L_0_inst : LUT6 generic map(INIT => "0000000001000100111011000000000000001101010000001100111100001000") port map( O =>C_48_S_1_L_0_out, I0 =>  inp_feat(33), I1 =>  inp_feat(22), I2 =>  inp_feat(469), I3 =>  inp_feat(253), I4 =>  inp_feat(289), I5 =>  inp_feat(13)); 
C_48_S_1_L_1_inst : LUT6 generic map(INIT => "0000100100000100000000011000110101101111001001011111011100011101") port map( O =>C_48_S_1_L_1_out, I0 =>  inp_feat(317), I1 =>  inp_feat(493), I2 =>  inp_feat(51), I3 =>  inp_feat(357), I4 =>  inp_feat(208), I5 =>  inp_feat(328)); 
C_48_S_1_L_2_inst : LUT6 generic map(INIT => "0001000000010000101100100001000010110111000110001111001101010011") port map( O =>C_48_S_1_L_2_out, I0 =>  inp_feat(246), I1 =>  inp_feat(469), I2 =>  inp_feat(354), I3 =>  inp_feat(197), I4 =>  inp_feat(385), I5 =>  inp_feat(13)); 
C_48_S_1_L_3_inst : LUT6 generic map(INIT => "0010000001110010100010100001000000000000000000000000000000010000") port map( O =>C_48_S_1_L_3_out, I0 =>  inp_feat(289), I1 =>  inp_feat(139), I2 =>  inp_feat(91), I3 =>  inp_feat(54), I4 =>  inp_feat(154), I5 =>  inp_feat(128)); 
C_48_S_1_L_4_inst : LUT6 generic map(INIT => "1111000101100001101001111000001100000000000000000000000000000001") port map( O =>C_48_S_1_L_4_out, I0 =>  inp_feat(115), I1 =>  inp_feat(375), I2 =>  inp_feat(288), I3 =>  inp_feat(192), I4 =>  inp_feat(368), I5 =>  inp_feat(128)); 
C_48_S_1_L_5_inst : LUT6 generic map(INIT => "0000100010100000000000000000100010110000111010000000000000000000") port map( O =>C_48_S_1_L_5_out, I0 =>  inp_feat(76), I1 =>  inp_feat(445), I2 =>  inp_feat(406), I3 =>  inp_feat(469), I4 =>  inp_feat(59), I5 =>  inp_feat(147)); 
C_48_S_2_L_0_inst : LUT6 generic map(INIT => "0000000000000010010001000110110111000100000001001100110011001101") port map( O =>C_48_S_2_L_0_out, I0 =>  inp_feat(413), I1 =>  inp_feat(189), I2 =>  inp_feat(33), I3 =>  inp_feat(380), I4 =>  inp_feat(51), I5 =>  inp_feat(328)); 
C_48_S_2_L_1_inst : LUT6 generic map(INIT => "0100000000010000000100001001000010110001111101000011000101110000") port map( O =>C_48_S_2_L_1_out, I0 =>  inp_feat(13), I1 =>  inp_feat(482), I2 =>  inp_feat(270), I3 =>  inp_feat(318), I4 =>  inp_feat(432), I5 =>  inp_feat(51)); 
C_48_S_2_L_2_inst : LUT6 generic map(INIT => "0000100101011111000001110001011111111111001101110011000101110111") port map( O =>C_48_S_2_L_2_out, I0 =>  inp_feat(48), I1 =>  inp_feat(183), I2 =>  inp_feat(249), I3 =>  inp_feat(81), I4 =>  inp_feat(509), I5 =>  inp_feat(448)); 
C_48_S_2_L_3_inst : LUT6 generic map(INIT => "0001000000110000000100101110000000000000110100000010110111011100") port map( O =>C_48_S_2_L_3_out, I0 =>  inp_feat(493), I1 =>  inp_feat(447), I2 =>  inp_feat(291), I3 =>  inp_feat(432), I4 =>  inp_feat(429), I5 =>  inp_feat(154)); 
C_48_S_2_L_4_inst : LUT6 generic map(INIT => "1001001011001001100011011100111100000000001000000000000000001110") port map( O =>C_48_S_2_L_4_out, I0 =>  inp_feat(415), I1 =>  inp_feat(383), I2 =>  inp_feat(89), I3 =>  inp_feat(263), I4 =>  inp_feat(378), I5 =>  inp_feat(389)); 
C_48_S_2_L_5_inst : LUT6 generic map(INIT => "0000010101110011000000000001000111010011001101010000010000000001") port map( O =>C_48_S_2_L_5_out, I0 =>  inp_feat(51), I1 =>  inp_feat(451), I2 =>  inp_feat(246), I3 =>  inp_feat(308), I4 =>  inp_feat(335), I5 =>  inp_feat(380)); 
C_48_S_3_L_0_inst : LUT6 generic map(INIT => "0001010000000100000001110111111110101101000001110111011101111111") port map( O =>C_48_S_3_L_0_out, I0 =>  inp_feat(139), I1 =>  inp_feat(378), I2 =>  inp_feat(413), I3 =>  inp_feat(418), I4 =>  inp_feat(66), I5 =>  inp_feat(208)); 
C_48_S_3_L_1_inst : LUT6 generic map(INIT => "0111000000010000110100000001100000000000000000000000000000000000") port map( O =>C_48_S_3_L_1_out, I0 =>  inp_feat(380), I1 =>  inp_feat(4), I2 =>  inp_feat(410), I3 =>  inp_feat(78), I4 =>  inp_feat(149), I5 =>  inp_feat(239)); 
C_48_S_3_L_2_inst : LUT6 generic map(INIT => "0001011100011111000101111101011100000011110101111010101100001111") port map( O =>C_48_S_3_L_2_out, I0 =>  inp_feat(81), I1 =>  inp_feat(453), I2 =>  inp_feat(183), I3 =>  inp_feat(149), I4 =>  inp_feat(429), I5 =>  inp_feat(375)); 
C_48_S_3_L_3_inst : LUT6 generic map(INIT => "1010110101010101000000000000001100000000000000000000000000000000") port map( O =>C_48_S_3_L_3_out, I0 =>  inp_feat(436), I1 =>  inp_feat(192), I2 =>  inp_feat(445), I3 =>  inp_feat(368), I4 =>  inp_feat(128), I5 =>  inp_feat(239)); 
C_48_S_3_L_4_inst : LUT6 generic map(INIT => "0010101011001000001101100000000110000010000010100000000010000001") port map( O =>C_48_S_3_L_4_out, I0 =>  inp_feat(296), I1 =>  inp_feat(151), I2 =>  inp_feat(51), I3 =>  inp_feat(33), I4 =>  inp_feat(160), I5 =>  inp_feat(343)); 
C_48_S_3_L_5_inst : LUT6 generic map(INIT => "0001001000000001000000000000000010010000111111110000000010101111") port map( O =>C_48_S_3_L_5_out, I0 =>  inp_feat(73), I1 =>  inp_feat(401), I2 =>  inp_feat(244), I3 =>  inp_feat(26), I4 =>  inp_feat(39), I5 =>  inp_feat(470)); 
C_48_S_4_L_0_inst : LUT6 generic map(INIT => "0101010100000101000000110000000111011111000101110000110111000111") port map( O =>C_48_S_4_L_0_out, I0 =>  inp_feat(81), I1 =>  inp_feat(89), I2 =>  inp_feat(183), I3 =>  inp_feat(254), I4 =>  inp_feat(332), I5 =>  inp_feat(208)); 
C_48_S_4_L_1_inst : LUT6 generic map(INIT => "0100000100001000011100010000000000000000000000000000000000000000") port map( O =>C_48_S_4_L_1_out, I0 =>  inp_feat(13), I1 =>  inp_feat(378), I2 =>  inp_feat(167), I3 =>  inp_feat(59), I4 =>  inp_feat(391), I5 =>  inp_feat(266)); 
C_48_S_4_L_2_inst : LUT6 generic map(INIT => "0101101101001111000000010100101100000000001111110100000000000001") port map( O =>C_48_S_4_L_2_out, I0 =>  inp_feat(378), I1 =>  inp_feat(183), I2 =>  inp_feat(469), I3 =>  inp_feat(317), I4 =>  inp_feat(372), I5 =>  inp_feat(236)); 
C_48_S_4_L_3_inst : LUT6 generic map(INIT => "1011111100000100000100111000000000000000000000000000000010000000") port map( O =>C_48_S_4_L_3_out, I0 =>  inp_feat(309), I1 =>  inp_feat(147), I2 =>  inp_feat(257), I3 =>  inp_feat(24), I4 =>  inp_feat(169), I5 =>  inp_feat(85)); 
C_48_S_4_L_4_inst : LUT6 generic map(INIT => "0101001000000010000100001000000001010100000000001100000000000000") port map( O =>C_48_S_4_L_4_out, I0 =>  inp_feat(380), I1 =>  inp_feat(359), I2 =>  inp_feat(140), I3 =>  inp_feat(60), I4 =>  inp_feat(372), I5 =>  inp_feat(236)); 
C_48_S_4_L_5_inst : LUT6 generic map(INIT => "1100011001110001000000001110101000000000000000000000000000000000") port map( O =>C_48_S_4_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(290), I2 =>  inp_feat(408), I3 =>  inp_feat(470), I4 =>  inp_feat(39), I5 =>  inp_feat(239)); 
C_48_S_5_L_0_inst : LUT6 generic map(INIT => "0011001000001010100000011010101000110000000000000010101100101110") port map( O =>C_48_S_5_L_0_out, I0 =>  inp_feat(339), I1 =>  inp_feat(215), I2 =>  inp_feat(250), I3 =>  inp_feat(91), I4 =>  inp_feat(366), I5 =>  inp_feat(77)); 
C_48_S_5_L_1_inst : LUT6 generic map(INIT => "0110000000000000000100000000001011110010111101100000000011100000") port map( O =>C_48_S_5_L_1_out, I0 =>  inp_feat(308), I1 =>  inp_feat(69), I2 =>  inp_feat(253), I3 =>  inp_feat(469), I4 =>  inp_feat(379), I5 =>  inp_feat(230)); 
C_48_S_5_L_2_inst : LUT6 generic map(INIT => "1001111101101111000000010100101100000000001111110100000000000001") port map( O =>C_48_S_5_L_2_out, I0 =>  inp_feat(378), I1 =>  inp_feat(183), I2 =>  inp_feat(469), I3 =>  inp_feat(317), I4 =>  inp_feat(372), I5 =>  inp_feat(236)); 
C_48_S_5_L_3_inst : LUT6 generic map(INIT => "0101111111100110000000111111011100000101000001010000010111000000") port map( O =>C_48_S_5_L_3_out, I0 =>  inp_feat(448), I1 =>  inp_feat(492), I2 =>  inp_feat(33), I3 =>  inp_feat(502), I4 =>  inp_feat(415), I5 =>  inp_feat(306)); 
C_48_S_5_L_4_inst : LUT6 generic map(INIT => "1001101100000100100100010000100100001000000000010000000000000000") port map( O =>C_48_S_5_L_4_out, I0 =>  inp_feat(210), I1 =>  inp_feat(407), I2 =>  inp_feat(429), I3 =>  inp_feat(383), I4 =>  inp_feat(420), I5 =>  inp_feat(199)); 
C_48_S_5_L_5_inst : LUT6 generic map(INIT => "0001010100000000000001000010000000000010000010010000000010000000") port map( O =>C_48_S_5_L_5_out, I0 =>  inp_feat(183), I1 =>  inp_feat(289), I2 =>  inp_feat(285), I3 =>  inp_feat(300), I4 =>  inp_feat(236), I5 =>  inp_feat(181)); 
C_49_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111100111111101110100011111110111111001110000011000000") port map( O =>C_49_S_0_L_0_out, I0 =>  inp_feat(151), I1 =>  inp_feat(183), I2 =>  inp_feat(246), I3 =>  inp_feat(378), I4 =>  inp_feat(317), I5 =>  inp_feat(469)); 
C_49_S_0_L_1_inst : LUT6 generic map(INIT => "1111101011010100111011111000100000000101000000001110101010000000") port map( O =>C_49_S_0_L_1_out, I0 =>  inp_feat(497), I1 =>  inp_feat(373), I2 =>  inp_feat(257), I3 =>  inp_feat(249), I4 =>  inp_feat(312), I5 =>  inp_feat(413)); 
C_49_S_0_L_2_inst : LUT6 generic map(INIT => "0000000011101101111111111110100011101110111011101110101010101010") port map( O =>C_49_S_0_L_2_out, I0 =>  inp_feat(438), I1 =>  inp_feat(493), I2 =>  inp_feat(378), I3 =>  inp_feat(503), I4 =>  inp_feat(52), I5 =>  inp_feat(420)); 
C_49_S_0_L_3_inst : LUT6 generic map(INIT => "1111111011111111001110111011011111101010111110100011001011111110") port map( O =>C_49_S_0_L_3_out, I0 =>  inp_feat(113), I1 =>  inp_feat(224), I2 =>  inp_feat(305), I3 =>  inp_feat(237), I4 =>  inp_feat(131), I5 =>  inp_feat(11)); 
C_49_S_0_L_4_inst : LUT6 generic map(INIT => "1111111111111111011100111111111100100011111100100111001111111011") port map( O =>C_49_S_0_L_4_out, I0 =>  inp_feat(411), I1 =>  inp_feat(94), I2 =>  inp_feat(348), I3 =>  inp_feat(323), I4 =>  inp_feat(435), I5 =>  inp_feat(352)); 
C_49_S_0_L_5_inst : LUT6 generic map(INIT => "1010110111111110000011001111100011111111111111111111111111111111") port map( O =>C_49_S_0_L_5_out, I0 =>  inp_feat(43), I1 =>  inp_feat(485), I2 =>  inp_feat(332), I3 =>  inp_feat(407), I4 =>  inp_feat(378), I5 =>  inp_feat(387)); 
C_49_S_1_L_0_inst : LUT6 generic map(INIT => "1110111111101110111000101110100000001100101011000000010010101000") port map( O =>C_49_S_1_L_0_out, I0 =>  inp_feat(328), I1 =>  inp_feat(81), I2 =>  inp_feat(72), I3 =>  inp_feat(312), I4 =>  inp_feat(445), I5 =>  inp_feat(413)); 
C_49_S_1_L_1_inst : LUT6 generic map(INIT => "1110001000000000111111101100100011111000111110101110100000001000") port map( O =>C_49_S_1_L_1_out, I0 =>  inp_feat(317), I1 =>  inp_feat(246), I2 =>  inp_feat(470), I3 =>  inp_feat(13), I4 =>  inp_feat(276), I5 =>  inp_feat(420)); 
C_49_S_1_L_2_inst : LUT6 generic map(INIT => "1111111100111110111111101010110000111110001011101111110011001100") port map( O =>C_49_S_1_L_2_out, I0 =>  inp_feat(130), I1 =>  inp_feat(39), I2 =>  inp_feat(224), I3 =>  inp_feat(230), I4 =>  inp_feat(190), I5 =>  inp_feat(147)); 
C_49_S_1_L_3_inst : LUT6 generic map(INIT => "0111011001110011111111111111001111101011110010001110100010000000") port map( O =>C_49_S_1_L_3_out, I0 =>  inp_feat(287), I1 =>  inp_feat(436), I2 =>  inp_feat(51), I3 =>  inp_feat(380), I4 =>  inp_feat(152), I5 =>  inp_feat(342)); 
C_49_S_1_L_4_inst : LUT6 generic map(INIT => "1100111011111110110001001110111001000000111100101000010011100000") port map( O =>C_49_S_1_L_4_out, I0 =>  inp_feat(469), I1 =>  inp_feat(51), I2 =>  inp_feat(352), I3 =>  inp_feat(130), I4 =>  inp_feat(476), I5 =>  inp_feat(378)); 
C_49_S_1_L_5_inst : LUT6 generic map(INIT => "1010101011011110111111001111100011101010111000100100111111111000") port map( O =>C_49_S_1_L_5_out, I0 =>  inp_feat(508), I1 =>  inp_feat(11), I2 =>  inp_feat(299), I3 =>  inp_feat(466), I4 =>  inp_feat(233), I5 =>  inp_feat(125)); 
C_49_S_2_L_0_inst : LUT6 generic map(INIT => "1000101001001101111110101111110011111111111110101111111010101000") port map( O =>C_49_S_2_L_0_out, I0 =>  inp_feat(156), I1 =>  inp_feat(317), I2 =>  inp_feat(125), I3 =>  inp_feat(208), I4 =>  inp_feat(127), I5 =>  inp_feat(454)); 
C_49_S_2_L_1_inst : LUT6 generic map(INIT => "1111111111111111100011101111111000101111111110110000101110100000") port map( O =>C_49_S_2_L_1_out, I0 =>  inp_feat(43), I1 =>  inp_feat(199), I2 =>  inp_feat(503), I3 =>  inp_feat(458), I4 =>  inp_feat(476), I5 =>  inp_feat(328)); 
C_49_S_2_L_2_inst : LUT6 generic map(INIT => "1111111110111001111111001111100000011101111101011100110000010000") port map( O =>C_49_S_2_L_2_out, I0 =>  inp_feat(185), I1 =>  inp_feat(204), I2 =>  inp_feat(487), I3 =>  inp_feat(305), I4 =>  inp_feat(379), I5 =>  inp_feat(469)); 
C_49_S_2_L_3_inst : LUT6 generic map(INIT => "1110100011111000111010111111111000000000001001101111111111101111") port map( O =>C_49_S_2_L_3_out, I0 =>  inp_feat(226), I1 =>  inp_feat(180), I2 =>  inp_feat(44), I3 =>  inp_feat(330), I4 =>  inp_feat(163), I5 =>  inp_feat(508)); 
C_49_S_2_L_4_inst : LUT6 generic map(INIT => "1101110111111110111111111110011100011110001010101111111111111111") port map( O =>C_49_S_2_L_4_out, I0 =>  inp_feat(485), I1 =>  inp_feat(178), I2 =>  inp_feat(356), I3 =>  inp_feat(291), I4 =>  inp_feat(420), I5 =>  inp_feat(289)); 
C_49_S_2_L_5_inst : LUT6 generic map(INIT => "0001000000100010111011001111011111111110111111101010000010000000") port map( O =>C_49_S_2_L_5_out, I0 =>  inp_feat(456), I1 =>  inp_feat(501), I2 =>  inp_feat(357), I3 =>  inp_feat(411), I4 =>  inp_feat(86), I5 =>  inp_feat(379)); 
C_49_S_3_L_0_inst : LUT6 generic map(INIT => "1110101011111100011110001111111011111101111110001110011001101100") port map( O =>C_49_S_3_L_0_out, I0 =>  inp_feat(84), I1 =>  inp_feat(418), I2 =>  inp_feat(33), I3 =>  inp_feat(365), I4 =>  inp_feat(330), I5 =>  inp_feat(94)); 
C_49_S_3_L_1_inst : LUT6 generic map(INIT => "0101100101000001111110010101110111111111111111111100111111100001") port map( O =>C_49_S_3_L_1_out, I0 =>  inp_feat(266), I1 =>  inp_feat(180), I2 =>  inp_feat(16), I3 =>  inp_feat(151), I4 =>  inp_feat(390), I5 =>  inp_feat(163)); 
C_49_S_3_L_2_inst : LUT6 generic map(INIT => "1110101001010000101110001100100011111111111111111010101000001000") port map( O =>C_49_S_3_L_2_out, I0 =>  inp_feat(81), I1 =>  inp_feat(51), I2 =>  inp_feat(249), I3 =>  inp_feat(508), I4 =>  inp_feat(183), I5 =>  inp_feat(454)); 
C_49_S_3_L_3_inst : LUT6 generic map(INIT => "0011001010101000101110001100000011111111111111111110111011101000") port map( O =>C_49_S_3_L_3_out, I0 =>  inp_feat(151), I1 =>  inp_feat(81), I2 =>  inp_feat(317), I3 =>  inp_feat(249), I4 =>  inp_feat(50), I5 =>  inp_feat(78)); 
C_49_S_3_L_4_inst : LUT6 generic map(INIT => "0110110010111100111010101111100011111101111011001111110000110000") port map( O =>C_49_S_3_L_4_out, I0 =>  inp_feat(249), I1 =>  inp_feat(373), I2 =>  inp_feat(51), I3 =>  inp_feat(508), I4 =>  inp_feat(183), I5 =>  inp_feat(454)); 
C_49_S_3_L_5_inst : LUT6 generic map(INIT => "1101010111011101111101011100111011001000001110001000101011110001") port map( O =>C_49_S_3_L_5_out, I0 =>  inp_feat(199), I1 =>  inp_feat(263), I2 =>  inp_feat(493), I3 =>  inp_feat(357), I4 =>  inp_feat(37), I5 =>  inp_feat(378)); 
C_49_S_4_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111110111101100000100000011101111010110111110") port map( O =>C_49_S_4_L_0_out, I0 =>  inp_feat(471), I1 =>  inp_feat(510), I2 =>  inp_feat(357), I3 =>  inp_feat(53), I4 =>  inp_feat(94), I5 =>  inp_feat(11)); 
C_49_S_4_L_1_inst : LUT6 generic map(INIT => "1110011101110011011101110110001101111011111100011111111110000000") port map( O =>C_49_S_4_L_1_out, I0 =>  inp_feat(480), I1 =>  inp_feat(420), I2 =>  inp_feat(289), I3 =>  inp_feat(33), I4 =>  inp_feat(492), I5 =>  inp_feat(401)); 
C_49_S_4_L_2_inst : LUT6 generic map(INIT => "1011011000110010001111111011001011111111101100100010001100100000") port map( O =>C_49_S_4_L_2_out, I0 =>  inp_feat(328), I1 =>  inp_feat(15), I2 =>  inp_feat(373), I3 =>  inp_feat(51), I4 =>  inp_feat(248), I5 =>  inp_feat(486)); 
C_49_S_4_L_3_inst : LUT6 generic map(INIT => "1000001111111000111111100110000001100101101000001011111010000000") port map( O =>C_49_S_4_L_3_out, I0 =>  inp_feat(125), I1 =>  inp_feat(390), I2 =>  inp_feat(208), I3 =>  inp_feat(382), I4 =>  inp_feat(39), I5 =>  inp_feat(328)); 
C_49_S_4_L_4_inst : LUT6 generic map(INIT => "1111000111110111101001111111111100001101101100111111111111110011") port map( O =>C_49_S_4_L_4_out, I0 =>  inp_feat(283), I1 =>  inp_feat(123), I2 =>  inp_feat(89), I3 =>  inp_feat(253), I4 =>  inp_feat(234), I5 =>  inp_feat(251)); 
C_49_S_4_L_5_inst : LUT6 generic map(INIT => "0100110100001001110101001111010111111111111111111100110010001000") port map( O =>C_49_S_4_L_5_out, I0 =>  inp_feat(190), I1 =>  inp_feat(317), I2 =>  inp_feat(249), I3 =>  inp_feat(411), I4 =>  inp_feat(183), I5 =>  inp_feat(454)); 
C_49_S_5_L_0_inst : LUT6 generic map(INIT => "1100111111110101110111001101001111111111111111101111111000111110") port map( O =>C_49_S_5_L_0_out, I0 =>  inp_feat(1), I1 =>  inp_feat(250), I2 =>  inp_feat(485), I3 =>  inp_feat(332), I4 =>  inp_feat(126), I5 =>  inp_feat(407)); 
C_49_S_5_L_1_inst : LUT6 generic map(INIT => "0111100111101101011111011110111111111101111111101111111111001111") port map( O =>C_49_S_5_L_1_out, I0 =>  inp_feat(95), I1 =>  inp_feat(485), I2 =>  inp_feat(401), I3 =>  inp_feat(332), I4 =>  inp_feat(43), I5 =>  inp_feat(407)); 
C_49_S_5_L_2_inst : LUT6 generic map(INIT => "1100001010110111111010001101110000101011010011000010100011111000") port map( O =>C_49_S_5_L_2_out, I0 =>  inp_feat(151), I1 =>  inp_feat(380), I2 =>  inp_feat(328), I3 =>  inp_feat(218), I4 =>  inp_feat(61), I5 =>  inp_feat(156)); 
C_49_S_5_L_3_inst : LUT6 generic map(INIT => "1000101011111000111001001111101011111111111110111000100000000000") port map( O =>C_49_S_5_L_3_out, I0 =>  inp_feat(51), I1 =>  inp_feat(451), I2 =>  inp_feat(470), I3 =>  inp_feat(276), I4 =>  inp_feat(111), I5 =>  inp_feat(22)); 
C_49_S_5_L_4_inst : LUT6 generic map(INIT => "1110011101010001111111110111110111111111001111101111001111111111") port map( O =>C_49_S_5_L_4_out, I0 =>  inp_feat(218), I1 =>  inp_feat(127), I2 =>  inp_feat(61), I3 =>  inp_feat(306), I4 =>  inp_feat(262), I5 =>  inp_feat(219)); 
C_49_S_5_L_5_inst : LUT6 generic map(INIT => "0110101011111110111011101100001000100010001110101110111100000000") port map( O =>C_49_S_5_L_5_out, I0 =>  inp_feat(249), I1 =>  inp_feat(372), I2 =>  inp_feat(276), I3 =>  inp_feat(111), I4 =>  inp_feat(22), I5 =>  inp_feat(451)); 
C_50_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111101110111111101110100011111110111000001110100000000000") port map( O =>C_50_S_0_L_0_out, I0 =>  inp_feat(378), I1 =>  inp_feat(183), I2 =>  inp_feat(249), I3 =>  inp_feat(246), I4 =>  inp_feat(84), I5 =>  inp_feat(469)); 
C_50_S_0_L_1_inst : LUT6 generic map(INIT => "0000011011001000001111111111111011111110111010000100001011100000") port map( O =>C_50_S_0_L_1_out, I0 =>  inp_feat(378), I1 =>  inp_feat(317), I2 =>  inp_feat(476), I3 =>  inp_feat(89), I4 =>  inp_feat(101), I5 =>  inp_feat(436)); 
C_50_S_0_L_2_inst : LUT6 generic map(INIT => "1011111000100000011110111110100011111110111110001111111111011100") port map( O =>C_50_S_0_L_2_out, I0 =>  inp_feat(131), I1 =>  inp_feat(451), I2 =>  inp_feat(69), I3 =>  inp_feat(373), I4 =>  inp_feat(190), I5 =>  inp_feat(18)); 
C_50_S_0_L_3_inst : LUT6 generic map(INIT => "0010100000000000101110001011110111111100111011100111111111111000") port map( O =>C_50_S_0_L_3_out, I0 =>  inp_feat(178), I1 =>  inp_feat(108), I2 =>  inp_feat(172), I3 =>  inp_feat(100), I4 =>  inp_feat(190), I5 =>  inp_feat(127)); 
C_50_S_0_L_4_inst : LUT6 generic map(INIT => "0111111001101000011111111010101011111110111010001111110011001000") port map( O =>C_50_S_0_L_4_out, I0 =>  inp_feat(246), I1 =>  inp_feat(378), I2 =>  inp_feat(149), I3 =>  inp_feat(375), I4 =>  inp_feat(301), I5 =>  inp_feat(45)); 
C_50_S_0_L_5_inst : LUT6 generic map(INIT => "1111111111101110111011101000100001101100111001001110000010000000") port map( O =>C_50_S_0_L_5_out, I0 =>  inp_feat(328), I1 =>  inp_feat(51), I2 =>  inp_feat(66), I3 =>  inp_feat(317), I4 =>  inp_feat(469), I5 =>  inp_feat(476)); 
C_50_S_1_L_0_inst : LUT6 generic map(INIT => "0000011011001000001111111111111011111110111010000100001011100000") port map( O =>C_50_S_1_L_0_out, I0 =>  inp_feat(378), I1 =>  inp_feat(317), I2 =>  inp_feat(476), I3 =>  inp_feat(89), I4 =>  inp_feat(101), I5 =>  inp_feat(436)); 
C_50_S_1_L_1_inst : LUT6 generic map(INIT => "1011111000100000011110111110100011111110111110001111111111011100") port map( O =>C_50_S_1_L_1_out, I0 =>  inp_feat(131), I1 =>  inp_feat(451), I2 =>  inp_feat(69), I3 =>  inp_feat(373), I4 =>  inp_feat(190), I5 =>  inp_feat(18)); 
C_50_S_1_L_2_inst : LUT6 generic map(INIT => "0010100000000000101110001011110111111100111011100111111111111000") port map( O =>C_50_S_1_L_2_out, I0 =>  inp_feat(178), I1 =>  inp_feat(108), I2 =>  inp_feat(172), I3 =>  inp_feat(100), I4 =>  inp_feat(190), I5 =>  inp_feat(127)); 
C_50_S_1_L_3_inst : LUT6 generic map(INIT => "0111111001101000011111111010101011111110111010001111110011001000") port map( O =>C_50_S_1_L_3_out, I0 =>  inp_feat(246), I1 =>  inp_feat(378), I2 =>  inp_feat(149), I3 =>  inp_feat(375), I4 =>  inp_feat(301), I5 =>  inp_feat(45)); 
C_50_S_1_L_4_inst : LUT6 generic map(INIT => "1111111111101110111011101000100001101100111001001110000010000000") port map( O =>C_50_S_1_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(51), I2 =>  inp_feat(66), I3 =>  inp_feat(317), I4 =>  inp_feat(469), I5 =>  inp_feat(476)); 
C_50_S_1_L_5_inst : LUT6 generic map(INIT => "0111111011111000000010110000000011111100111110000001000010110000") port map( O =>C_50_S_1_L_5_out, I0 =>  inp_feat(246), I1 =>  inp_feat(378), I2 =>  inp_feat(183), I3 =>  inp_feat(81), I4 =>  inp_feat(305), I5 =>  inp_feat(296)); 
C_50_S_2_L_0_inst : LUT6 generic map(INIT => "0001111011011110111111101100100011111110110000001110000000000000") port map( O =>C_50_S_2_L_0_out, I0 =>  inp_feat(435), I1 =>  inp_feat(246), I2 =>  inp_feat(13), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_2_L_1_inst : LUT6 generic map(INIT => "1101111111101110111111101110100011111111100010001110000010000000") port map( O =>C_50_S_2_L_1_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_2_L_2_inst : LUT6 generic map(INIT => "0000110101101010011010100110101010111111100010001100000000000000") port map( O =>C_50_S_2_L_2_out, I0 =>  inp_feat(373), I1 =>  inp_feat(13), I2 =>  inp_feat(289), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_2_L_3_inst : LUT6 generic map(INIT => "1111111111101110111111101110100011111010100011001110000010000000") port map( O =>C_50_S_2_L_3_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_2_L_4_inst : LUT6 generic map(INIT => "0111111101001110011111101100100011111010100010001110000010000000") port map( O =>C_50_S_2_L_4_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_2_L_5_inst : LUT6 generic map(INIT => "1011111100101110111111101110100001011110100001001110000010000000") port map( O =>C_50_S_2_L_5_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_3_L_0_inst : LUT6 generic map(INIT => "1111010001101100011011001110110011111110111010001110000010100000") port map( O =>C_50_S_3_L_0_out, I0 =>  inp_feat(51), I1 =>  inp_feat(373), I2 =>  inp_feat(13), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_3_L_1_inst : LUT6 generic map(INIT => "0001101111101110111111101100100011111010100010001110000010000000") port map( O =>C_50_S_3_L_1_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_3_L_2_inst : LUT6 generic map(INIT => "1101110100101110111111101110100011111111100011001110000010000000") port map( O =>C_50_S_3_L_2_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_3_L_3_inst : LUT6 generic map(INIT => "0011001111001110011111101100100011111010100010001110000010000000") port map( O =>C_50_S_3_L_3_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_3_L_4_inst : LUT6 generic map(INIT => "1100111001111010011010100110101001111110100010001110000000000000") port map( O =>C_50_S_3_L_4_out, I0 =>  inp_feat(413), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_3_L_5_inst : LUT6 generic map(INIT => "0011000111000010111111101100100001011010100001001110000010000000") port map( O =>C_50_S_3_L_5_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_4_L_0_inst : LUT6 generic map(INIT => "0001101001101100111011100110110011011110111010001110000010100000") port map( O =>C_50_S_4_L_0_out, I0 =>  inp_feat(51), I1 =>  inp_feat(373), I2 =>  inp_feat(13), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_4_L_1_inst : LUT6 generic map(INIT => "1101111110101110111111101110100011111010100011001110000010000000") port map( O =>C_50_S_4_L_1_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_4_L_2_inst : LUT6 generic map(INIT => "0011101111101110010111101100100011111010100010001110000010000000") port map( O =>C_50_S_4_L_2_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_4_L_3_inst : LUT6 generic map(INIT => "0100111000111010011010100110101011111110100010001110000000000000") port map( O =>C_50_S_4_L_3_out, I0 =>  inp_feat(413), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_4_L_4_inst : LUT6 generic map(INIT => "1101000101000010111101101100100001111011100001001110000010000000") port map( O =>C_50_S_4_L_4_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_4_L_5_inst : LUT6 generic map(INIT => "0111011111011110011010101110100001100110100010001110000000000000") port map( O =>C_50_S_4_L_5_out, I0 =>  inp_feat(413), I1 =>  inp_feat(131), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_5_L_0_inst : LUT6 generic map(INIT => "1101111110100110111111101110100011111110100010001110000010000000") port map( O =>C_50_S_5_L_0_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_5_L_1_inst : LUT6 generic map(INIT => "0010111011111010011010100100101011111110100010001110000000000000") port map( O =>C_50_S_5_L_1_out, I0 =>  inp_feat(413), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_5_L_2_inst : LUT6 generic map(INIT => "1101100100100010110101101110100001011010100011001110000010000000") port map( O =>C_50_S_5_L_2_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_5_L_3_inst : LUT6 generic map(INIT => "0110011011001010011010100101101011111110100010001110000000000000") port map( O =>C_50_S_5_L_3_out, I0 =>  inp_feat(413), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_5_L_4_inst : LUT6 generic map(INIT => "1010001001011010111110100110101001111000010010001100000010000000") port map( O =>C_50_S_5_L_4_out, I0 =>  inp_feat(435), I1 =>  inp_feat(317), I2 =>  inp_feat(13), I3 =>  inp_feat(246), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_50_S_5_L_5_inst : LUT6 generic map(INIT => "0111110100101110010101100100100001110010100001001110000010000000") port map( O =>C_50_S_5_L_5_out, I0 =>  inp_feat(51), I1 =>  inp_feat(246), I2 =>  inp_feat(147), I3 =>  inp_feat(317), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_51_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111110111011101110100011111110111111001111000011100000") port map( O =>C_51_S_0_L_0_out, I0 =>  inp_feat(183), I1 =>  inp_feat(378), I2 =>  inp_feat(317), I3 =>  inp_feat(51), I4 =>  inp_feat(246), I5 =>  inp_feat(469)); 
C_51_S_0_L_1_inst : LUT6 generic map(INIT => "1101111011011110000101001111110100000010010110100010000011110000") port map( O =>C_51_S_0_L_1_out, I0 =>  inp_feat(281), I1 =>  inp_feat(304), I2 =>  inp_feat(413), I3 =>  inp_feat(426), I4 =>  inp_feat(81), I5 =>  inp_feat(249)); 
C_51_S_0_L_2_inst : LUT6 generic map(INIT => "1011111111111101000011001111111000100111111101110000001011101100") port map( O =>C_51_S_0_L_2_out, I0 =>  inp_feat(33), I1 =>  inp_feat(183), I2 =>  inp_feat(180), I3 =>  inp_feat(312), I4 =>  inp_feat(151), I5 =>  inp_feat(343)); 
C_51_S_0_L_3_inst : LUT6 generic map(INIT => "1110111100111110011111100000100000001000001011000110100000001000") port map( O =>C_51_S_0_L_3_out, I0 =>  inp_feat(78), I1 =>  inp_feat(335), I2 =>  inp_feat(253), I3 =>  inp_feat(51), I4 =>  inp_feat(373), I5 =>  inp_feat(11)); 
C_51_S_0_L_4_inst : LUT6 generic map(INIT => "1101100101001110010111100101110011111111111111101111000011001101") port map( O =>C_51_S_0_L_4_out, I0 =>  inp_feat(305), I1 =>  inp_feat(50), I2 =>  inp_feat(221), I3 =>  inp_feat(446), I4 =>  inp_feat(263), I5 =>  inp_feat(272)); 
C_51_S_0_L_5_inst : LUT6 generic map(INIT => "1011000010000000101100101100100010111100100000000010010000000000") port map( O =>C_51_S_0_L_5_out, I0 =>  inp_feat(147), I1 =>  inp_feat(469), I2 =>  inp_feat(246), I3 =>  inp_feat(413), I4 =>  inp_feat(28), I5 =>  inp_feat(117)); 
C_51_S_1_L_0_inst : LUT6 generic map(INIT => "1101111011011110000101001111110100000010010110100010000011110000") port map( O =>C_51_S_1_L_0_out, I0 =>  inp_feat(281), I1 =>  inp_feat(304), I2 =>  inp_feat(413), I3 =>  inp_feat(426), I4 =>  inp_feat(81), I5 =>  inp_feat(249)); 
C_51_S_1_L_1_inst : LUT6 generic map(INIT => "1011111111111101000011001111111000100111111101110000001011101100") port map( O =>C_51_S_1_L_1_out, I0 =>  inp_feat(33), I1 =>  inp_feat(183), I2 =>  inp_feat(180), I3 =>  inp_feat(312), I4 =>  inp_feat(151), I5 =>  inp_feat(343)); 
C_51_S_1_L_2_inst : LUT6 generic map(INIT => "1110111100111110011111100000100000001000001011000110100000001000") port map( O =>C_51_S_1_L_2_out, I0 =>  inp_feat(78), I1 =>  inp_feat(335), I2 =>  inp_feat(253), I3 =>  inp_feat(51), I4 =>  inp_feat(373), I5 =>  inp_feat(11)); 
C_51_S_1_L_3_inst : LUT6 generic map(INIT => "1101100101001110010111100101110011111111111111101111000011001101") port map( O =>C_51_S_1_L_3_out, I0 =>  inp_feat(305), I1 =>  inp_feat(50), I2 =>  inp_feat(221), I3 =>  inp_feat(446), I4 =>  inp_feat(263), I5 =>  inp_feat(272)); 
C_51_S_1_L_4_inst : LUT6 generic map(INIT => "1011000010000000101100101100100010111100100000000010010000000000") port map( O =>C_51_S_1_L_4_out, I0 =>  inp_feat(147), I1 =>  inp_feat(469), I2 =>  inp_feat(246), I3 =>  inp_feat(413), I4 =>  inp_feat(28), I5 =>  inp_feat(117)); 
C_51_S_1_L_5_inst : LUT6 generic map(INIT => "1011000111110111101111110001110100010101111111011111010000000011") port map( O =>C_51_S_1_L_5_out, I0 =>  inp_feat(59), I1 =>  inp_feat(283), I2 =>  inp_feat(418), I3 =>  inp_feat(248), I4 =>  inp_feat(187), I5 =>  inp_feat(163)); 
C_51_S_2_L_0_inst : LUT6 generic map(INIT => "0111000010000000011001101111001011111111111111101111111111001000") port map( O =>C_51_S_2_L_0_out, I0 =>  inp_feat(13), I1 =>  inp_feat(435), I2 =>  inp_feat(413), I3 =>  inp_feat(195), I4 =>  inp_feat(180), I5 =>  inp_feat(312)); 
C_51_S_2_L_1_inst : LUT6 generic map(INIT => "1000111011111010011000111111000011111011111111111101001111111111") port map( O =>C_51_S_2_L_1_out, I0 =>  inp_feat(296), I1 =>  inp_feat(180), I2 =>  inp_feat(176), I3 =>  inp_feat(464), I4 =>  inp_feat(258), I5 =>  inp_feat(232)); 
C_51_S_2_L_2_inst : LUT6 generic map(INIT => "1011101111111010001100111111111000110010110011000000000011000100") port map( O =>C_51_S_2_L_2_out, I0 =>  inp_feat(183), I1 =>  inp_feat(237), I2 =>  inp_feat(329), I3 =>  inp_feat(253), I4 =>  inp_feat(51), I5 =>  inp_feat(373)); 
C_51_S_2_L_3_inst : LUT6 generic map(INIT => "0111110100101011010011100111011111111111111111111111111100111010") port map( O =>C_51_S_2_L_3_out, I0 =>  inp_feat(375), I1 =>  inp_feat(112), I2 =>  inp_feat(306), I3 =>  inp_feat(215), I4 =>  inp_feat(242), I5 =>  inp_feat(181)); 
C_51_S_2_L_4_inst : LUT6 generic map(INIT => "1100111011110000111111000111110100100010101000001111110111111111") port map( O =>C_51_S_2_L_4_out, I0 =>  inp_feat(51), I1 =>  inp_feat(33), I2 =>  inp_feat(413), I3 =>  inp_feat(230), I4 =>  inp_feat(323), I5 =>  inp_feat(469)); 
C_51_S_2_L_5_inst : LUT6 generic map(INIT => "1011101101011110100011100111101010110110011010001110111000001000") port map( O =>C_51_S_2_L_5_out, I0 =>  inp_feat(7), I1 =>  inp_feat(426), I2 =>  inp_feat(419), I3 =>  inp_feat(246), I4 =>  inp_feat(348), I5 =>  inp_feat(163)); 
C_51_S_3_L_0_inst : LUT6 generic map(INIT => "0001010101101110001000001110110011111111111011101111001101001010") port map( O =>C_51_S_3_L_0_out, I0 =>  inp_feat(148), I1 =>  inp_feat(491), I2 =>  inp_feat(60), I3 =>  inp_feat(72), I4 =>  inp_feat(180), I5 =>  inp_feat(312)); 
C_51_S_3_L_1_inst : LUT6 generic map(INIT => "1111010111101100111111101110110011111111000011000101000011010100") port map( O =>C_51_S_3_L_1_out, I0 =>  inp_feat(510), I1 =>  inp_feat(446), I2 =>  inp_feat(105), I3 =>  inp_feat(389), I4 =>  inp_feat(8), I5 =>  inp_feat(226)); 
C_51_S_3_L_2_inst : LUT6 generic map(INIT => "1000000100010100111111000110100011111010111111101111111100001110") port map( O =>C_51_S_3_L_2_out, I0 =>  inp_feat(160), I1 =>  inp_feat(249), I2 =>  inp_feat(81), I3 =>  inp_feat(222), I4 =>  inp_feat(351), I5 =>  inp_feat(59)); 
C_51_S_3_L_3_inst : LUT6 generic map(INIT => "0000011111010101100000011001111011110111110111111111111100101111") port map( O =>C_51_S_3_L_3_out, I0 =>  inp_feat(415), I1 =>  inp_feat(180), I2 =>  inp_feat(238), I3 =>  inp_feat(484), I4 =>  inp_feat(38), I5 =>  inp_feat(232)); 
C_51_S_3_L_4_inst : LUT6 generic map(INIT => "1010111100101110111111111110101000001110000011111111111001011100") port map( O =>C_51_S_3_L_4_out, I0 =>  inp_feat(77), I1 =>  inp_feat(96), I2 =>  inp_feat(312), I3 =>  inp_feat(289), I4 =>  inp_feat(142), I5 =>  inp_feat(38)); 
C_51_S_3_L_5_inst : LUT6 generic map(INIT => "0101100010111110000111001111000011111000111110100110000011110000") port map( O =>C_51_S_3_L_5_out, I0 =>  inp_feat(492), I1 =>  inp_feat(84), I2 =>  inp_feat(51), I3 =>  inp_feat(306), I4 =>  inp_feat(365), I5 =>  inp_feat(486)); 
C_51_S_4_L_0_inst : LUT6 generic map(INIT => "0101111111111111110110011000110000110111010111111111111110111100") port map( O =>C_51_S_4_L_0_out, I0 =>  inp_feat(216), I1 =>  inp_feat(176), I2 =>  inp_feat(138), I3 =>  inp_feat(494), I4 =>  inp_feat(379), I5 =>  inp_feat(434)); 
C_51_S_4_L_1_inst : LUT6 generic map(INIT => "1100001010100000111001111111111111111011111001101111111110001111") port map( O =>C_51_S_4_L_1_out, I0 =>  inp_feat(378), I1 =>  inp_feat(113), I2 =>  inp_feat(470), I3 =>  inp_feat(446), I4 =>  inp_feat(399), I5 =>  inp_feat(279)); 
C_51_S_4_L_2_inst : LUT6 generic map(INIT => "1011001011001110111111000111110000110010000111101110110010000000") port map( O =>C_51_S_4_L_2_out, I0 =>  inp_feat(435), I1 =>  inp_feat(334), I2 =>  inp_feat(42), I3 =>  inp_feat(127), I4 =>  inp_feat(101), I5 =>  inp_feat(258)); 
C_51_S_4_L_3_inst : LUT6 generic map(INIT => "1111110100001110111011101100101010001100110001101000000001001010") port map( O =>C_51_S_4_L_3_out, I0 =>  inp_feat(478), I1 =>  inp_feat(51), I2 =>  inp_feat(46), I3 =>  inp_feat(99), I4 =>  inp_feat(57), I5 =>  inp_feat(50)); 
C_51_S_4_L_4_inst : LUT6 generic map(INIT => "0000101011000001110111111111111111111111111010001111111011111000") port map( O =>C_51_S_4_L_4_out, I0 =>  inp_feat(264), I1 =>  inp_feat(230), I2 =>  inp_feat(459), I3 =>  inp_feat(79), I4 =>  inp_feat(232), I5 =>  inp_feat(114)); 
C_51_S_4_L_5_inst : LUT6 generic map(INIT => "1010111110101111111111111101101000000011111110001110110010000000") port map( O =>C_51_S_4_L_5_out, I0 =>  inp_feat(258), I1 =>  inp_feat(288), I2 =>  inp_feat(191), I3 =>  inp_feat(383), I4 =>  inp_feat(306), I5 =>  inp_feat(163)); 
C_51_S_5_L_0_inst : LUT6 generic map(INIT => "1111111111111111011011111111111000011000111110011111110011001000") port map( O =>C_51_S_5_L_0_out, I0 =>  inp_feat(479), I1 =>  inp_feat(128), I2 =>  inp_feat(405), I3 =>  inp_feat(282), I4 =>  inp_feat(434), I5 =>  inp_feat(296)); 
C_51_S_5_L_1_inst : LUT6 generic map(INIT => "0010000011111100010110001111100011111000111111111111111010001101") port map( O =>C_51_S_5_L_1_out, I0 =>  inp_feat(208), I1 =>  inp_feat(249), I2 =>  inp_feat(438), I3 =>  inp_feat(234), I4 =>  inp_feat(176), I5 =>  inp_feat(15)); 
C_51_S_5_L_2_inst : LUT6 generic map(INIT => "1110110011110110010100101111011100101010111010001110111011101110") port map( O =>C_51_S_5_L_2_out, I0 =>  inp_feat(51), I1 =>  inp_feat(380), I2 =>  inp_feat(289), I3 =>  inp_feat(279), I4 =>  inp_feat(207), I5 =>  inp_feat(453)); 
C_51_S_5_L_3_inst : LUT6 generic map(INIT => "0001001110000010001100111011000111111111111100111111000011000001") port map( O =>C_51_S_5_L_3_out, I0 =>  inp_feat(289), I1 =>  inp_feat(136), I2 =>  inp_feat(131), I3 =>  inp_feat(385), I4 =>  inp_feat(469), I5 =>  inp_feat(326)); 
C_51_S_5_L_4_inst : LUT6 generic map(INIT => "1000111010101010000011001101101000011111111011101111111011101101") port map( O =>C_51_S_5_L_4_out, I0 =>  inp_feat(328), I1 =>  inp_feat(33), I2 =>  inp_feat(64), I3 =>  inp_feat(305), I4 =>  inp_feat(93), I5 =>  inp_feat(0)); 
C_51_S_5_L_5_inst : LUT6 generic map(INIT => "1111101010101010110010001110001000000100110010001110110011000000") port map( O =>C_51_S_5_L_5_out, I0 =>  inp_feat(81), I1 =>  inp_feat(289), I2 =>  inp_feat(328), I3 =>  inp_feat(89), I4 =>  inp_feat(423), I5 =>  inp_feat(476)); 
C_52_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000011000000000001011100010001000101110000000101111111") port map( O =>C_52_S_0_L_0_out, I0 =>  inp_feat(317), I1 =>  inp_feat(378), I2 =>  inp_feat(328), I3 =>  inp_feat(51), I4 =>  inp_feat(84), I5 =>  inp_feat(469)); 
C_52_S_0_L_1_inst : LUT6 generic map(INIT => "0000000100100011110001011110001110000111001111111000000000010111") port map( O =>C_52_S_0_L_1_out, I0 =>  inp_feat(50), I1 =>  inp_feat(317), I2 =>  inp_feat(289), I3 =>  inp_feat(246), I4 =>  inp_feat(321), I5 =>  inp_feat(470)); 
C_52_S_0_L_2_inst : LUT6 generic map(INIT => "1010100011101110111011001111111100000000110011001100111011100000") port map( O =>C_52_S_0_L_2_out, I0 =>  inp_feat(182), I1 =>  inp_feat(413), I2 =>  inp_feat(422), I3 =>  inp_feat(218), I4 =>  inp_feat(163), I5 =>  inp_feat(37)); 
C_52_S_0_L_3_inst : LUT6 generic map(INIT => "0001000001010001010111001111000111011100000010000010000001010000") port map( O =>C_52_S_0_L_3_out, I0 =>  inp_feat(413), I1 =>  inp_feat(208), I2 =>  inp_feat(182), I3 =>  inp_feat(469), I4 =>  inp_feat(380), I5 =>  inp_feat(227)); 
C_52_S_0_L_4_inst : LUT6 generic map(INIT => "1100001011000110000000101100000000000010000000000000001001000100") port map( O =>C_52_S_0_L_4_out, I0 =>  inp_feat(90), I1 =>  inp_feat(246), I2 =>  inp_feat(413), I3 =>  inp_feat(488), I4 =>  inp_feat(78), I5 =>  inp_feat(461)); 
C_52_S_0_L_5_inst : LUT6 generic map(INIT => "0000001001110111000100001011100100101000011111010001100011111001") port map( O =>C_52_S_0_L_5_out, I0 =>  inp_feat(151), I1 =>  inp_feat(50), I2 =>  inp_feat(509), I3 =>  inp_feat(13), I4 =>  inp_feat(389), I5 =>  inp_feat(171)); 
C_52_S_1_L_0_inst : LUT6 generic map(INIT => "0000000000010101101000001001010110000001000101111000000000010111") port map( O =>C_52_S_1_L_0_out, I0 =>  inp_feat(317), I1 =>  inp_feat(51), I2 =>  inp_feat(289), I3 =>  inp_feat(246), I4 =>  inp_feat(321), I5 =>  inp_feat(470)); 
C_52_S_1_L_1_inst : LUT6 generic map(INIT => "1011001111000100111101111100100001010101000000001101011110000000") port map( O =>C_52_S_1_L_1_out, I0 =>  inp_feat(289), I1 =>  inp_feat(469), I2 =>  inp_feat(418), I3 =>  inp_feat(22), I4 =>  inp_feat(171), I5 =>  inp_feat(37)); 
C_52_S_1_L_2_inst : LUT6 generic map(INIT => "0000000001010101000100011010001100111100001110110101111100111111") port map( O =>C_52_S_1_L_2_out, I0 =>  inp_feat(435), I1 =>  inp_feat(51), I2 =>  inp_feat(373), I3 =>  inp_feat(131), I4 =>  inp_feat(230), I5 =>  inp_feat(289)); 
C_52_S_1_L_3_inst : LUT6 generic map(INIT => "1101000000000111110110111010111100100000001000110000001100011111") port map( O =>C_52_S_1_L_3_out, I0 =>  inp_feat(453), I1 =>  inp_feat(154), I2 =>  inp_feat(350), I3 =>  inp_feat(503), I4 =>  inp_feat(204), I5 =>  inp_feat(480)); 
C_52_S_1_L_4_inst : LUT6 generic map(INIT => "0101100001010001010101001111000000000000000000000000000000010001") port map( O =>C_52_S_1_L_4_out, I0 =>  inp_feat(103), I1 =>  inp_feat(90), I2 =>  inp_feat(413), I3 =>  inp_feat(488), I4 =>  inp_feat(78), I5 =>  inp_feat(461)); 
C_52_S_1_L_5_inst : LUT6 generic map(INIT => "1011111011101111101001011101110110110010001000000000000000001101") port map( O =>C_52_S_1_L_5_out, I0 =>  inp_feat(378), I1 =>  inp_feat(293), I2 =>  inp_feat(447), I3 =>  inp_feat(89), I4 =>  inp_feat(11), I5 =>  inp_feat(182)); 
C_52_S_2_L_0_inst : LUT6 generic map(INIT => "0101100100100010000110111010101111010001000000100011000100001011") port map( O =>C_52_S_2_L_0_out, I0 =>  inp_feat(420), I1 =>  inp_feat(13), I2 =>  inp_feat(378), I3 =>  inp_feat(246), I4 =>  inp_feat(469), I5 =>  inp_feat(218)); 
C_52_S_2_L_1_inst : LUT6 generic map(INIT => "1110110011000000010101011111011101100000110100000011000111110001") port map( O =>C_52_S_2_L_1_out, I0 =>  inp_feat(131), I1 =>  inp_feat(230), I2 =>  inp_feat(222), I3 =>  inp_feat(50), I4 =>  inp_feat(139), I5 =>  inp_feat(117)); 
C_52_S_2_L_2_inst : LUT6 generic map(INIT => "0000010100111111000001110011111110101001100110010001111101111111") port map( O =>C_52_S_2_L_2_out, I0 =>  inp_feat(151), I1 =>  inp_feat(413), I2 =>  inp_feat(131), I3 =>  inp_feat(246), I4 =>  inp_feat(139), I5 =>  inp_feat(385)); 
C_52_S_2_L_3_inst : LUT6 generic map(INIT => "1001011100011111100000000000100011011011110111111010100010000000") port map( O =>C_52_S_2_L_3_out, I0 =>  inp_feat(435), I1 =>  inp_feat(249), I2 =>  inp_feat(469), I3 =>  inp_feat(380), I4 =>  inp_feat(68), I5 =>  inp_feat(412)); 
C_52_S_2_L_4_inst : LUT6 generic map(INIT => "0000100100010111000000011011011100001101000111110000011111111111") port map( O =>C_52_S_2_L_4_out, I0 =>  inp_feat(435), I1 =>  inp_feat(413), I2 =>  inp_feat(13), I3 =>  inp_feat(246), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_52_S_2_L_5_inst : LUT6 generic map(INIT => "0011000000001001000001000000100011111111101100100101000000001000") port map( O =>C_52_S_2_L_5_out, I0 =>  inp_feat(111), I1 =>  inp_feat(190), I2 =>  inp_feat(483), I3 =>  inp_feat(372), I4 =>  inp_feat(324), I5 =>  inp_feat(163)); 
C_52_S_3_L_0_inst : LUT6 generic map(INIT => "1110000000010010011000111100000111001101000001111001111101111111") port map( O =>C_52_S_3_L_0_out, I0 =>  inp_feat(373), I1 =>  inp_feat(378), I2 =>  inp_feat(413), I3 =>  inp_feat(380), I4 =>  inp_feat(131), I5 =>  inp_feat(51)); 
C_52_S_3_L_1_inst : LUT6 generic map(INIT => "1100000011100101010010010001011100101100010111010011111111111111") port map( O =>C_52_S_3_L_1_out, I0 =>  inp_feat(317), I1 =>  inp_feat(208), I2 =>  inp_feat(13), I3 =>  inp_feat(246), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_52_S_3_L_2_inst : LUT6 generic map(INIT => "0000001011110000111100001010000001010000110101001001010100101111") port map( O =>C_52_S_3_L_2_out, I0 =>  inp_feat(401), I1 =>  inp_feat(307), I2 =>  inp_feat(46), I3 =>  inp_feat(502), I4 =>  inp_feat(163), I5 =>  inp_feat(287)); 
C_52_S_3_L_3_inst : LUT6 generic map(INIT => "0010011010100011100010101011001101000110001010110010111110111111") port map( O =>C_52_S_3_L_3_out, I0 =>  inp_feat(389), I1 =>  inp_feat(413), I2 =>  inp_feat(13), I3 =>  inp_feat(246), I4 =>  inp_feat(380), I5 =>  inp_feat(469)); 
C_52_S_3_L_4_inst : LUT6 generic map(INIT => "0110100000001100011101000000000011111000000000001111001001110000") port map( O =>C_52_S_3_L_4_out, I0 =>  inp_feat(227), I1 =>  inp_feat(405), I2 =>  inp_feat(493), I3 =>  inp_feat(376), I4 =>  inp_feat(175), I5 =>  inp_feat(220)); 
C_52_S_3_L_5_inst : LUT6 generic map(INIT => "0111011110110001000100111000000111011001110100111101001100010001") port map( O =>C_52_S_3_L_5_out, I0 =>  inp_feat(81), I1 =>  inp_feat(13), I2 =>  inp_feat(195), I3 =>  inp_feat(31), I4 =>  inp_feat(330), I5 =>  inp_feat(456)); 
C_52_S_4_L_0_inst : LUT6 generic map(INIT => "1100101001011000011100000110000000101011001100010111110011110101") port map( O =>C_52_S_4_L_0_out, I0 =>  inp_feat(469), I1 =>  inp_feat(482), I2 =>  inp_feat(22), I3 =>  inp_feat(413), I4 =>  inp_feat(246), I5 =>  inp_feat(51)); 
C_52_S_4_L_1_inst : LUT6 generic map(INIT => "0100111000111010001000111011001001100000101010100011101011111111") port map( O =>C_52_S_4_L_1_out, I0 =>  inp_feat(234), I1 =>  inp_feat(434), I2 =>  inp_feat(385), I3 =>  inp_feat(413), I4 =>  inp_feat(246), I5 =>  inp_feat(51)); 
C_52_S_4_L_2_inst : LUT6 generic map(INIT => "1000001100000001110100111111111110100011101000111001111111111111") port map( O =>C_52_S_4_L_2_out, I0 =>  inp_feat(13), I1 =>  inp_feat(183), I2 =>  inp_feat(151), I3 =>  inp_feat(413), I4 =>  inp_feat(246), I5 =>  inp_feat(352)); 
C_52_S_4_L_3_inst : LUT6 generic map(INIT => "1110010000001100101100000011000000010100000000001011001001000000") port map( O =>C_52_S_4_L_3_out, I0 =>  inp_feat(13), I1 =>  inp_feat(55), I2 =>  inp_feat(249), I3 =>  inp_feat(376), I4 =>  inp_feat(220), I5 =>  inp_feat(330)); 
C_52_S_4_L_4_inst : LUT6 generic map(INIT => "0000000101000010010110110001000110101001000001111101110101111111") port map( O =>C_52_S_4_L_4_out, I0 =>  inp_feat(317), I1 =>  inp_feat(378), I2 =>  inp_feat(435), I3 =>  inp_feat(380), I4 =>  inp_feat(131), I5 =>  inp_feat(51)); 
C_52_S_4_L_5_inst : LUT6 generic map(INIT => "1000110011000111111011100010101100000000010010111010010100010111") port map( O =>C_52_S_4_L_5_out, I0 =>  inp_feat(235), I1 =>  inp_feat(106), I2 =>  inp_feat(369), I3 =>  inp_feat(17), I4 =>  inp_feat(141), I5 =>  inp_feat(192)); 
C_52_S_5_L_0_inst : LUT6 generic map(INIT => "1101101100101111110110001000110000000010000011001000100000001110") port map( O =>C_52_S_5_L_0_out, I0 =>  inp_feat(89), I1 =>  inp_feat(322), I2 =>  inp_feat(336), I3 =>  inp_feat(17), I4 =>  inp_feat(162), I5 =>  inp_feat(472)); 
C_52_S_5_L_1_inst : LUT6 generic map(INIT => "0101111101001001101011001000000000000001000000010100110010001101") port map( O =>C_52_S_5_L_1_out, I0 =>  inp_feat(490), I1 =>  inp_feat(436), I2 =>  inp_feat(191), I3 =>  inp_feat(502), I4 =>  inp_feat(163), I5 =>  inp_feat(287)); 
C_52_S_5_L_2_inst : LUT6 generic map(INIT => "0100010100000010000101000000110010000100111111110001110011001110") port map( O =>C_52_S_5_L_2_out, I0 =>  inp_feat(404), I1 =>  inp_feat(221), I2 =>  inp_feat(317), I3 =>  inp_feat(183), I4 =>  inp_feat(373), I5 =>  inp_feat(98)); 
C_52_S_5_L_3_inst : LUT6 generic map(INIT => "1100010111000001100101110111111110000000010000010000000100000001") port map( O =>C_52_S_5_L_3_out, I0 =>  inp_feat(435), I1 =>  inp_feat(183), I2 =>  inp_feat(451), I3 =>  inp_feat(50), I4 =>  inp_feat(139), I5 =>  inp_feat(201)); 
C_52_S_5_L_4_inst : LUT6 generic map(INIT => "0000101000000000010110010010000010010000000111011101100001000000") port map( O =>C_52_S_5_L_4_out, I0 =>  inp_feat(183), I1 =>  inp_feat(135), I2 =>  inp_feat(338), I3 =>  inp_feat(221), I4 =>  inp_feat(378), I5 =>  inp_feat(434)); 
C_52_S_5_L_5_inst : LUT6 generic map(INIT => "1000110111111111000101000101110111011111001111110100110000111111") port map( O =>C_52_S_5_L_5_out, I0 =>  inp_feat(166), I1 =>  inp_feat(343), I2 =>  inp_feat(175), I3 =>  inp_feat(412), I4 =>  inp_feat(38), I5 =>  inp_feat(220)); 
C_53_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000011000000010001011100010001000101110000000101111111") port map( O =>C_53_S_0_L_0_out, I0 =>  inp_feat(317), I1 =>  inp_feat(378), I2 =>  inp_feat(328), I3 =>  inp_feat(51), I4 =>  inp_feat(84), I5 =>  inp_feat(469)); 
C_53_S_0_L_1_inst : LUT6 generic map(INIT => "1000110110011101000000010000110000000000000001010000000000001100") port map( O =>C_53_S_0_L_1_out, I0 =>  inp_feat(471), I1 =>  inp_feat(221), I2 =>  inp_feat(413), I3 =>  inp_feat(375), I4 =>  inp_feat(332), I5 =>  inp_feat(419)); 
C_53_S_0_L_2_inst : LUT6 generic map(INIT => "1111100011001000110100001110110000000000100000000000000000100000") port map( O =>C_53_S_0_L_2_out, I0 =>  inp_feat(32), I1 =>  inp_feat(291), I2 =>  inp_feat(436), I3 =>  inp_feat(434), I4 =>  inp_feat(147), I5 =>  inp_feat(488)); 
C_53_S_0_L_3_inst : LUT6 generic map(INIT => "0000001111010011000100011101000100000000000000010000010000000011") port map( O =>C_53_S_0_L_3_out, I0 =>  inp_feat(394), I1 =>  inp_feat(160), I2 =>  inp_feat(68), I3 =>  inp_feat(330), I4 =>  inp_feat(49), I5 =>  inp_feat(189)); 
C_53_S_0_L_4_inst : LUT6 generic map(INIT => "0101101011111000011100011111110000000000100100000000000001100000") port map( O =>C_53_S_0_L_4_out, I0 =>  inp_feat(469), I1 =>  inp_feat(456), I2 =>  inp_feat(393), I3 =>  inp_feat(413), I4 =>  inp_feat(51), I5 =>  inp_feat(455)); 
C_53_S_0_L_5_inst : LUT6 generic map(INIT => "1010111100011101111000101101000000000000000000101110000000000000") port map( O =>C_53_S_0_L_5_out, I0 =>  inp_feat(403), I1 =>  inp_feat(413), I2 =>  inp_feat(472), I3 =>  inp_feat(232), I4 =>  inp_feat(246), I5 =>  inp_feat(483)); 
C_53_S_1_L_0_inst : LUT6 generic map(INIT => "1000110110011101000000010000110000000000000001010000000000001100") port map( O =>C_53_S_1_L_0_out, I0 =>  inp_feat(471), I1 =>  inp_feat(221), I2 =>  inp_feat(413), I3 =>  inp_feat(375), I4 =>  inp_feat(332), I5 =>  inp_feat(419)); 
C_53_S_1_L_1_inst : LUT6 generic map(INIT => "1111100011001000110100001110110000000000100000000000000000100000") port map( O =>C_53_S_1_L_1_out, I0 =>  inp_feat(32), I1 =>  inp_feat(291), I2 =>  inp_feat(436), I3 =>  inp_feat(434), I4 =>  inp_feat(147), I5 =>  inp_feat(488)); 
C_53_S_1_L_2_inst : LUT6 generic map(INIT => "0000001111010011000100011101000100000000000000010000010000000011") port map( O =>C_53_S_1_L_2_out, I0 =>  inp_feat(394), I1 =>  inp_feat(160), I2 =>  inp_feat(68), I3 =>  inp_feat(330), I4 =>  inp_feat(49), I5 =>  inp_feat(189)); 
C_53_S_1_L_3_inst : LUT6 generic map(INIT => "0101101011111000011100011111110000000000100100000000000001100000") port map( O =>C_53_S_1_L_3_out, I0 =>  inp_feat(469), I1 =>  inp_feat(456), I2 =>  inp_feat(393), I3 =>  inp_feat(413), I4 =>  inp_feat(51), I5 =>  inp_feat(455)); 
C_53_S_1_L_4_inst : LUT6 generic map(INIT => "1010111100011101111000101101000000000000000000101110000000000000") port map( O =>C_53_S_1_L_4_out, I0 =>  inp_feat(403), I1 =>  inp_feat(413), I2 =>  inp_feat(472), I3 =>  inp_feat(232), I4 =>  inp_feat(246), I5 =>  inp_feat(483)); 
C_53_S_1_L_5_inst : LUT6 generic map(INIT => "1010001010101000101010101011000000010000000010000000000011100010") port map( O =>C_53_S_1_L_5_out, I0 =>  inp_feat(426), I1 =>  inp_feat(50), I2 =>  inp_feat(1), I3 =>  inp_feat(264), I4 =>  inp_feat(13), I5 =>  inp_feat(189)); 
C_53_S_2_L_0_inst : LUT6 generic map(INIT => "1101010111100001010101110001000000000100100111000001000000001000") port map( O =>C_53_S_2_L_0_out, I0 =>  inp_feat(246), I1 =>  inp_feat(151), I2 =>  inp_feat(138), I3 =>  inp_feat(481), I4 =>  inp_feat(391), I5 =>  inp_feat(455)); 
C_53_S_2_L_1_inst : LUT6 generic map(INIT => "0100110011010101001000000010000001000001110000000001000000000000") port map( O =>C_53_S_2_L_1_out, I0 =>  inp_feat(475), I1 =>  inp_feat(480), I2 =>  inp_feat(375), I3 =>  inp_feat(502), I4 =>  inp_feat(468), I5 =>  inp_feat(39)); 
C_53_S_2_L_2_inst : LUT6 generic map(INIT => "1111001100000001111000111000000001110010000100000000000000000000") port map( O =>C_53_S_2_L_2_out, I0 =>  inp_feat(434), I1 =>  inp_feat(413), I2 =>  inp_feat(375), I3 =>  inp_feat(502), I4 =>  inp_feat(468), I5 =>  inp_feat(39)); 
C_53_S_2_L_3_inst : LUT6 generic map(INIT => "1111000111110100001110000011001000110001000001000000000000000000") port map( O =>C_53_S_2_L_3_out, I0 =>  inp_feat(127), I1 =>  inp_feat(505), I2 =>  inp_feat(144), I3 =>  inp_feat(11), I4 =>  inp_feat(111), I5 =>  inp_feat(483)); 
C_53_S_2_L_4_inst : LUT6 generic map(INIT => "0000000000000100101101001100000000000000000000001111110000000001") port map( O =>C_53_S_2_L_4_out, I0 =>  inp_feat(263), I1 =>  inp_feat(224), I2 =>  inp_feat(319), I3 =>  inp_feat(316), I4 =>  inp_feat(200), I5 =>  inp_feat(15)); 
C_53_S_2_L_5_inst : LUT6 generic map(INIT => "1001111010001010101111010010001000000110000000100000000000001100") port map( O =>C_53_S_2_L_5_out, I0 =>  inp_feat(338), I1 =>  inp_feat(208), I2 =>  inp_feat(416), I3 =>  inp_feat(418), I4 =>  inp_feat(476), I5 =>  inp_feat(458)); 
C_53_S_3_L_0_inst : LUT6 generic map(INIT => "0010010100010000110011000000000000010001111000001100011100100000") port map( O =>C_53_S_3_L_0_out, I0 =>  inp_feat(218), I1 =>  inp_feat(298), I2 =>  inp_feat(101), I3 =>  inp_feat(70), I4 =>  inp_feat(505), I5 =>  inp_feat(290)); 
C_53_S_3_L_1_inst : LUT6 generic map(INIT => "1100111001101110101010000010100000000100000001001101000000000000") port map( O =>C_53_S_3_L_1_out, I0 =>  inp_feat(17), I1 =>  inp_feat(90), I2 =>  inp_feat(257), I3 =>  inp_feat(468), I4 =>  inp_feat(167), I5 =>  inp_feat(306)); 
C_53_S_3_L_2_inst : LUT6 generic map(INIT => "0010000101010001011000101100100010001000110100001010111100000000") port map( O =>C_53_S_3_L_2_out, I0 =>  inp_feat(23), I1 =>  inp_feat(192), I2 =>  inp_feat(476), I3 =>  inp_feat(232), I4 =>  inp_feat(470), I5 =>  inp_feat(50)); 
C_53_S_3_L_3_inst : LUT6 generic map(INIT => "0010001100001011001010010001000111010011011111111010000100010111") port map( O =>C_53_S_3_L_3_out, I0 =>  inp_feat(317), I1 =>  inp_feat(246), I2 =>  inp_feat(51), I3 =>  inp_feat(289), I4 =>  inp_feat(489), I5 =>  inp_feat(215)); 
C_53_S_3_L_4_inst : LUT6 generic map(INIT => "1111000011110001011111101101100001010001011100010101000011011000") port map( O =>C_53_S_3_L_4_out, I0 =>  inp_feat(486), I1 =>  inp_feat(141), I2 =>  inp_feat(441), I3 =>  inp_feat(487), I4 =>  inp_feat(54), I5 =>  inp_feat(29)); 
C_53_S_3_L_5_inst : LUT6 generic map(INIT => "1000100011000101011011011000110000000010010100000000000000001000") port map( O =>C_53_S_3_L_5_out, I0 =>  inp_feat(11), I1 =>  inp_feat(187), I2 =>  inp_feat(144), I3 =>  inp_feat(413), I4 =>  inp_feat(323), I5 =>  inp_feat(115)); 
C_53_S_4_L_0_inst : LUT6 generic map(INIT => "1000101010000110001100101010000010000000000000010000000000000010") port map( O =>C_53_S_4_L_0_out, I0 =>  inp_feat(111), I1 =>  inp_feat(231), I2 =>  inp_feat(250), I3 =>  inp_feat(200), I4 =>  inp_feat(503), I5 =>  inp_feat(290)); 
C_53_S_4_L_1_inst : LUT6 generic map(INIT => "0101000111110000011000000111000000110001001000101011000000101000") port map( O =>C_53_S_4_L_1_out, I0 =>  inp_feat(250), I1 =>  inp_feat(470), I2 =>  inp_feat(290), I3 =>  inp_feat(352), I4 =>  inp_feat(331), I5 =>  inp_feat(316)); 
C_53_S_4_L_2_inst : LUT6 generic map(INIT => "1111010110001001011001011000100001000001100100000000000000001000") port map( O =>C_53_S_4_L_2_out, I0 =>  inp_feat(205), I1 =>  inp_feat(224), I2 =>  inp_feat(136), I3 =>  inp_feat(460), I4 =>  inp_feat(296), I5 =>  inp_feat(316)); 
C_53_S_4_L_3_inst : LUT6 generic map(INIT => "1000100110001000001010001110111000000000000010000000100010001100") port map( O =>C_53_S_4_L_3_out, I0 =>  inp_feat(85), I1 =>  inp_feat(403), I2 =>  inp_feat(236), I3 =>  inp_feat(413), I4 =>  inp_feat(69), I5 =>  inp_feat(182)); 
C_53_S_4_L_4_inst : LUT6 generic map(INIT => "0001000000100000000110110110000000011011000000011111111100000011") port map( O =>C_53_S_4_L_4_out, I0 =>  inp_feat(209), I1 =>  inp_feat(413), I2 =>  inp_feat(482), I3 =>  inp_feat(253), I4 =>  inp_feat(435), I5 =>  inp_feat(69)); 
C_53_S_4_L_5_inst : LUT6 generic map(INIT => "1011111110110101110111000100000100010001110100000000000000110000") port map( O =>C_53_S_4_L_5_out, I0 =>  inp_feat(161), I1 =>  inp_feat(334), I2 =>  inp_feat(489), I3 =>  inp_feat(487), I4 =>  inp_feat(476), I5 =>  inp_feat(44)); 
C_53_S_5_L_0_inst : LUT6 generic map(INIT => "0000000010000010000100101001100010010010000000111100001101110000") port map( O =>C_53_S_5_L_0_out, I0 =>  inp_feat(199), I1 =>  inp_feat(133), I2 =>  inp_feat(154), I3 =>  inp_feat(174), I4 =>  inp_feat(383), I5 =>  inp_feat(200)); 
C_53_S_5_L_1_inst : LUT6 generic map(INIT => "1111001000001010111100000110001000000000000010001111001000100100") port map( O =>C_53_S_5_L_1_out, I0 =>  inp_feat(131), I1 =>  inp_feat(195), I2 =>  inp_feat(112), I3 =>  inp_feat(22), I4 =>  inp_feat(0), I5 =>  inp_feat(458)); 
C_53_S_5_L_2_inst : LUT6 generic map(INIT => "1010111010000001011011110000010000000000000100000101110100001100") port map( O =>C_53_S_5_L_2_out, I0 =>  inp_feat(283), I1 =>  inp_feat(489), I2 =>  inp_feat(472), I3 =>  inp_feat(92), I4 =>  inp_feat(161), I5 =>  inp_feat(182)); 
C_53_S_5_L_3_inst : LUT6 generic map(INIT => "0000000101001001110001001010000001010011001001101000010000000000") port map( O =>C_53_S_5_L_3_out, I0 =>  inp_feat(67), I1 =>  inp_feat(386), I2 =>  inp_feat(465), I3 =>  inp_feat(419), I4 =>  inp_feat(303), I5 =>  inp_feat(110)); 
C_53_S_5_L_4_inst : LUT6 generic map(INIT => "1000000010010100111110010010100000000000000000110111001110000000") port map( O =>C_53_S_5_L_4_out, I0 =>  inp_feat(164), I1 =>  inp_feat(106), I2 =>  inp_feat(475), I3 =>  inp_feat(480), I4 =>  inp_feat(136), I5 =>  inp_feat(115)); 
C_53_S_5_L_5_inst : LUT6 generic map(INIT => "0000010100000001001001000000110011011101010001000000110011111111") port map( O =>C_53_S_5_L_5_out, I0 =>  inp_feat(151), I1 =>  inp_feat(283), I2 =>  inp_feat(368), I3 =>  inp_feat(51), I4 =>  inp_feat(380), I5 =>  inp_feat(435)); 
C_54_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111101100111011001000100011111011111110101110100010000000") port map( O =>C_54_S_0_L_0_out, I0 =>  inp_feat(379), I1 =>  inp_feat(316), I2 =>  inp_feat(372), I3 =>  inp_feat(282), I4 =>  inp_feat(436), I5 =>  inp_feat(444)); 
C_54_S_0_L_1_inst : LUT6 generic map(INIT => "0011100001101000111011001100100011111111111100101110111100000001") port map( O =>C_54_S_0_L_1_out, I0 =>  inp_feat(104), I1 =>  inp_feat(312), I2 =>  inp_feat(432), I3 =>  inp_feat(282), I4 =>  inp_feat(183), I5 =>  inp_feat(438)); 
C_54_S_0_L_2_inst : LUT6 generic map(INIT => "0011111110101010011111111110100001011100100010001101100010000000") port map( O =>C_54_S_0_L_2_out, I0 =>  inp_feat(312), I1 =>  inp_feat(387), I2 =>  inp_feat(316), I3 =>  inp_feat(173), I4 =>  inp_feat(282), I5 =>  inp_feat(432)); 
C_54_S_0_L_3_inst : LUT6 generic map(INIT => "1110100001101010101010001100000011101110101010101110100010000000") port map( O =>C_54_S_0_L_3_out, I0 =>  inp_feat(170), I1 =>  inp_feat(312), I2 =>  inp_feat(372), I3 =>  inp_feat(266), I4 =>  inp_feat(15), I5 =>  inp_feat(386)); 
C_54_S_0_L_4_inst : LUT6 generic map(INIT => "0111111101111010011011001100000001111110011010001110000010000000") port map( O =>C_54_S_0_L_4_out, I0 =>  inp_feat(379), I1 =>  inp_feat(221), I2 =>  inp_feat(372), I3 =>  inp_feat(432), I4 =>  inp_feat(104), I5 =>  inp_feat(444)); 
C_54_S_0_L_5_inst : LUT6 generic map(INIT => "1111111010011010111111001100000001111110001010000110000010000000") port map( O =>C_54_S_0_L_5_out, I0 =>  inp_feat(379), I1 =>  inp_feat(221), I2 =>  inp_feat(372), I3 =>  inp_feat(432), I4 =>  inp_feat(104), I5 =>  inp_feat(444)); 
C_54_S_1_L_0_inst : LUT6 generic map(INIT => "0011100001101000111011001100100011111111111100101110111100000001") port map( O =>C_54_S_1_L_0_out, I0 =>  inp_feat(104), I1 =>  inp_feat(312), I2 =>  inp_feat(432), I3 =>  inp_feat(282), I4 =>  inp_feat(183), I5 =>  inp_feat(438)); 
C_54_S_1_L_1_inst : LUT6 generic map(INIT => "1101010110101110111101101010001000010000101110100101001010100000") port map( O =>C_54_S_1_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(28), I2 =>  inp_feat(383), I3 =>  inp_feat(316), I4 =>  inp_feat(270), I5 =>  inp_feat(92)); 
C_54_S_1_L_2_inst : LUT6 generic map(INIT => "0010111010101000001011001110000011111110111010000001100001000000") port map( O =>C_54_S_1_L_2_out, I0 =>  inp_feat(432), I1 =>  inp_feat(379), I2 =>  inp_feat(316), I3 =>  inp_feat(387), I4 =>  inp_feat(266), I5 =>  inp_feat(386)); 
C_54_S_1_L_3_inst : LUT6 generic map(INIT => "1011111111111011111111001110100001111011110001001100100000000000") port map( O =>C_54_S_1_L_3_out, I0 =>  inp_feat(282), I1 =>  inp_feat(221), I2 =>  inp_feat(257), I3 =>  inp_feat(170), I4 =>  inp_feat(173), I5 =>  inp_feat(312)); 
C_54_S_1_L_4_inst : LUT6 generic map(INIT => "0100000001001101100111000101000011101101111100001010001000010000") port map( O =>C_54_S_1_L_4_out, I0 =>  inp_feat(195), I1 =>  inp_feat(82), I2 =>  inp_feat(20), I3 =>  inp_feat(342), I4 =>  inp_feat(58), I5 =>  inp_feat(301)); 
C_54_S_1_L_5_inst : LUT6 generic map(INIT => "0101010011110000111110001000000011111101110100001111000000000000") port map( O =>C_54_S_1_L_5_out, I0 =>  inp_feat(139), I1 =>  inp_feat(74), I2 =>  inp_feat(312), I3 =>  inp_feat(270), I4 =>  inp_feat(332), I5 =>  inp_feat(77)); 
C_54_S_2_L_0_inst : LUT6 generic map(INIT => "0111110001111110011010001010100000111100010011000010000010001000") port map( O =>C_54_S_2_L_0_out, I0 =>  inp_feat(379), I1 =>  inp_feat(312), I2 =>  inp_feat(173), I3 =>  inp_feat(470), I4 =>  inp_feat(257), I5 =>  inp_feat(270)); 
C_54_S_2_L_1_inst : LUT6 generic map(INIT => "0101110011010000111011001010000011101111111111101110110011100000") port map( O =>C_54_S_2_L_1_out, I0 =>  inp_feat(143), I1 =>  inp_feat(58), I2 =>  inp_feat(462), I3 =>  inp_feat(0), I4 =>  inp_feat(8), I5 =>  inp_feat(261)); 
C_54_S_2_L_2_inst : LUT6 generic map(INIT => "1011100111101001111111111101111100101011010110110100111001011100") port map( O =>C_54_S_2_L_2_out, I0 =>  inp_feat(319), I1 =>  inp_feat(379), I2 =>  inp_feat(419), I3 =>  inp_feat(170), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_2_L_3_inst : LUT6 generic map(INIT => "0001110011100010011111100011000011110011111011101111100010000000") port map( O =>C_54_S_2_L_3_out, I0 =>  inp_feat(74), I1 =>  inp_feat(175), I2 =>  inp_feat(173), I3 =>  inp_feat(221), I4 =>  inp_feat(363), I5 =>  inp_feat(49)); 
C_54_S_2_L_4_inst : LUT6 generic map(INIT => "1011011110111100101110111011000000111011110100000001110000000000") port map( O =>C_54_S_2_L_4_out, I0 =>  inp_feat(72), I1 =>  inp_feat(292), I2 =>  inp_feat(436), I3 =>  inp_feat(316), I4 =>  inp_feat(312), I5 =>  inp_feat(248)); 
C_54_S_2_L_5_inst : LUT6 generic map(INIT => "0011111011111000110011001100100010111110111110001110000011000000") port map( O =>C_54_S_2_L_5_out, I0 =>  inp_feat(257), I1 =>  inp_feat(379), I2 =>  inp_feat(221), I3 =>  inp_feat(372), I4 =>  inp_feat(391), I5 =>  inp_feat(317)); 
C_54_S_3_L_0_inst : LUT6 generic map(INIT => "0110110111101111111001101000111001110110110010000010111100000000") port map( O =>C_54_S_3_L_0_out, I0 =>  inp_feat(418), I1 =>  inp_feat(312), I2 =>  inp_feat(165), I3 =>  inp_feat(316), I4 =>  inp_feat(379), I5 =>  inp_feat(266)); 
C_54_S_3_L_1_inst : LUT6 generic map(INIT => "1001100111011000001111101111100001001100000110100110110000000000") port map( O =>C_54_S_3_L_1_out, I0 =>  inp_feat(300), I1 =>  inp_feat(176), I2 =>  inp_feat(165), I3 =>  inp_feat(316), I4 =>  inp_feat(266), I5 =>  inp_feat(379)); 
C_54_S_3_L_2_inst : LUT6 generic map(INIT => "0011110111001011111110101010101001101110010010101100000000000000") port map( O =>C_54_S_3_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(76), I2 =>  inp_feat(368), I3 =>  inp_feat(316), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_3_L_3_inst : LUT6 generic map(INIT => "1111010011011101101111111101111101010111110100001101101101000000") port map( O =>C_54_S_3_L_3_out, I0 =>  inp_feat(215), I1 =>  inp_feat(316), I2 =>  inp_feat(454), I3 =>  inp_feat(173), I4 =>  inp_feat(282), I5 =>  inp_feat(432)); 
C_54_S_3_L_4_inst : LUT6 generic map(INIT => "0111110111111100111011001111110000011111111110000000000010100000") port map( O =>C_54_S_3_L_4_out, I0 =>  inp_feat(54), I1 =>  inp_feat(226), I2 =>  inp_feat(394), I3 =>  inp_feat(319), I4 =>  inp_feat(253), I5 =>  inp_feat(257)); 
C_54_S_3_L_5_inst : LUT6 generic map(INIT => "1111111101111111010110111010101000111110110010001100000000001000") port map( O =>C_54_S_3_L_5_out, I0 =>  inp_feat(221), I1 =>  inp_feat(170), I2 =>  inp_feat(368), I3 =>  inp_feat(316), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_4_L_0_inst : LUT6 generic map(INIT => "1111110011011110111100101110100010001110100011101100000000000000") port map( O =>C_54_S_4_L_0_out, I0 =>  inp_feat(316), I1 =>  inp_feat(432), I2 =>  inp_feat(334), I3 =>  inp_feat(253), I4 =>  inp_feat(257), I5 =>  inp_feat(270)); 
C_54_S_4_L_1_inst : LUT6 generic map(INIT => "0011111101111111110110111010101000011110010010001110000000001000") port map( O =>C_54_S_4_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(170), I2 =>  inp_feat(368), I3 =>  inp_feat(316), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_4_L_2_inst : LUT6 generic map(INIT => "1111111001101010111110100000000000011000010010001011100011000000") port map( O =>C_54_S_4_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(130), I2 =>  inp_feat(221), I3 =>  inp_feat(312), I4 =>  inp_feat(32), I5 =>  inp_feat(105)); 
C_54_S_4_L_3_inst : LUT6 generic map(INIT => "0010001000001010100000100110000011111010000000001111001001110000") port map( O =>C_54_S_4_L_3_out, I0 =>  inp_feat(274), I1 =>  inp_feat(169), I2 =>  inp_feat(248), I3 =>  inp_feat(170), I4 =>  inp_feat(312), I5 =>  inp_feat(10)); 
C_54_S_4_L_4_inst : LUT6 generic map(INIT => "1111001110011111101110111010101000111110010010001110000000001000") port map( O =>C_54_S_4_L_4_out, I0 =>  inp_feat(221), I1 =>  inp_feat(170), I2 =>  inp_feat(368), I3 =>  inp_feat(316), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_4_L_5_inst : LUT6 generic map(INIT => "0100001001101011000000010101111110101010101110000010001011101101") port map( O =>C_54_S_4_L_5_out, I0 =>  inp_feat(275), I1 =>  inp_feat(479), I2 =>  inp_feat(415), I3 =>  inp_feat(26), I4 =>  inp_feat(143), I5 =>  inp_feat(23)); 
C_54_S_5_L_0_inst : LUT6 generic map(INIT => "1101101011101110011111101110111001101000101000001110000010000000") port map( O =>C_54_S_5_L_0_out, I0 =>  inp_feat(170), I1 =>  inp_feat(257), I2 =>  inp_feat(363), I3 =>  inp_feat(282), I4 =>  inp_feat(173), I5 =>  inp_feat(221)); 
C_54_S_5_L_1_inst : LUT6 generic map(INIT => "1101001011010111101011001010111101100111001101110010111000000010") port map( O =>C_54_S_5_L_1_out, I0 =>  inp_feat(379), I1 =>  inp_feat(124), I2 =>  inp_feat(419), I3 =>  inp_feat(316), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_5_L_2_inst : LUT6 generic map(INIT => "0001001110111011000110111010101000111110010010001100000000001000") port map( O =>C_54_S_5_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(170), I2 =>  inp_feat(368), I3 =>  inp_feat(316), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_54_S_5_L_3_inst : LUT6 generic map(INIT => "0101111111011000110111001110100001011101100101000101010000000000") port map( O =>C_54_S_5_L_3_out, I0 =>  inp_feat(470), I1 =>  inp_feat(432), I2 =>  inp_feat(102), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_54_S_5_L_4_inst : LUT6 generic map(INIT => "1111110100000011101101111101111110110101010101110001111100010000") port map( O =>C_54_S_5_L_4_out, I0 =>  inp_feat(450), I1 =>  inp_feat(262), I2 =>  inp_feat(92), I3 =>  inp_feat(221), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_54_S_5_L_5_inst : LUT6 generic map(INIT => "0000101101001110110100010000110011101000111010001110010000000000") port map( O =>C_54_S_5_L_5_out, I0 =>  inp_feat(334), I1 =>  inp_feat(170), I2 =>  inp_feat(395), I3 =>  inp_feat(221), I4 =>  inp_feat(248), I5 =>  inp_feat(405)); 
C_55_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000000001001100000001000101110001111101111111") port map( O =>C_55_S_0_L_0_out, I0 =>  inp_feat(312), I1 =>  inp_feat(170), I2 =>  inp_feat(248), I3 =>  inp_feat(221), I4 =>  inp_feat(379), I5 =>  inp_feat(316)); 
C_55_S_0_L_1_inst : LUT6 generic map(INIT => "0001001000000000010111010000100011111111001000000000000000000000") port map( O =>C_55_S_0_L_1_out, I0 =>  inp_feat(432), I1 =>  inp_feat(157), I2 =>  inp_feat(351), I3 =>  inp_feat(11), I4 =>  inp_feat(204), I5 =>  inp_feat(173)); 
C_55_S_0_L_2_inst : LUT6 generic map(INIT => "0101111100000011111101010000001100000001000000000011000100000000") port map( O =>C_55_S_0_L_2_out, I0 =>  inp_feat(282), I1 =>  inp_feat(170), I2 =>  inp_feat(257), I3 =>  inp_feat(20), I4 =>  inp_feat(461), I5 =>  inp_feat(456)); 
C_55_S_0_L_3_inst : LUT6 generic map(INIT => "0101000100010001100111110100111100000000001100000010000100000111") port map( O =>C_55_S_0_L_3_out, I0 =>  inp_feat(266), I1 =>  inp_feat(493), I2 =>  inp_feat(157), I3 =>  inp_feat(311), I4 =>  inp_feat(180), I5 =>  inp_feat(11)); 
C_55_S_0_L_4_inst : LUT6 generic map(INIT => "0000001101010000000100111101001011011101000001010000000011000000") port map( O =>C_55_S_0_L_4_out, I0 =>  inp_feat(170), I1 =>  inp_feat(101), I2 =>  inp_feat(316), I3 =>  inp_feat(450), I4 =>  inp_feat(454), I5 =>  inp_feat(387)); 
C_55_S_0_L_5_inst : LUT6 generic map(INIT => "1001110000001000111101110000000000000000000000000111000000001000") port map( O =>C_55_S_0_L_5_out, I0 =>  inp_feat(311), I1 =>  inp_feat(187), I2 =>  inp_feat(139), I3 =>  inp_feat(169), I4 =>  inp_feat(121), I5 =>  inp_feat(71)); 
C_55_S_1_L_0_inst : LUT6 generic map(INIT => "0001001000000000010111010000100011111111001000000000000000000000") port map( O =>C_55_S_1_L_0_out, I0 =>  inp_feat(432), I1 =>  inp_feat(157), I2 =>  inp_feat(351), I3 =>  inp_feat(11), I4 =>  inp_feat(204), I5 =>  inp_feat(173)); 
C_55_S_1_L_1_inst : LUT6 generic map(INIT => "0101111100000011111101010000001100000001000000000011000100000000") port map( O =>C_55_S_1_L_1_out, I0 =>  inp_feat(282), I1 =>  inp_feat(170), I2 =>  inp_feat(257), I3 =>  inp_feat(20), I4 =>  inp_feat(461), I5 =>  inp_feat(456)); 
C_55_S_1_L_2_inst : LUT6 generic map(INIT => "0101000100010001100111110100111100000000001100000010000100000111") port map( O =>C_55_S_1_L_2_out, I0 =>  inp_feat(266), I1 =>  inp_feat(493), I2 =>  inp_feat(157), I3 =>  inp_feat(311), I4 =>  inp_feat(180), I5 =>  inp_feat(11)); 
C_55_S_1_L_3_inst : LUT6 generic map(INIT => "0000001101010000000100111101001011011101000001010000000011000000") port map( O =>C_55_S_1_L_3_out, I0 =>  inp_feat(170), I1 =>  inp_feat(101), I2 =>  inp_feat(316), I3 =>  inp_feat(450), I4 =>  inp_feat(454), I5 =>  inp_feat(387)); 
C_55_S_1_L_4_inst : LUT6 generic map(INIT => "1001110000001000111101110000000000000000000000000111000000001000") port map( O =>C_55_S_1_L_4_out, I0 =>  inp_feat(311), I1 =>  inp_feat(187), I2 =>  inp_feat(139), I3 =>  inp_feat(169), I4 =>  inp_feat(121), I5 =>  inp_feat(71)); 
C_55_S_1_L_5_inst : LUT6 generic map(INIT => "0010000000001101100001010000100000000000100000101100101000100000") port map( O =>C_55_S_1_L_5_out, I0 =>  inp_feat(26), I1 =>  inp_feat(22), I2 =>  inp_feat(342), I3 =>  inp_feat(191), I4 =>  inp_feat(296), I5 =>  inp_feat(506)); 
C_55_S_2_L_0_inst : LUT6 generic map(INIT => "1110011000000111100101110001111100000001000000010000000110011111") port map( O =>C_55_S_2_L_0_out, I0 =>  inp_feat(253), I1 =>  inp_feat(379), I2 =>  inp_feat(387), I3 =>  inp_feat(432), I4 =>  inp_feat(257), I5 =>  inp_feat(20)); 
C_55_S_2_L_1_inst : LUT6 generic map(INIT => "0011111100001111000101010000001100010111000001110000000010000001") port map( O =>C_55_S_2_L_1_out, I0 =>  inp_feat(379), I1 =>  inp_feat(248), I2 =>  inp_feat(387), I3 =>  inp_feat(2), I4 =>  inp_feat(508), I5 =>  inp_feat(230)); 
C_55_S_2_L_2_inst : LUT6 generic map(INIT => "0000010001001100000000000010110011111101011101000000001001100100") port map( O =>C_55_S_2_L_2_out, I0 =>  inp_feat(253), I1 =>  inp_feat(399), I2 =>  inp_feat(506), I3 =>  inp_feat(366), I4 =>  inp_feat(228), I5 =>  inp_feat(112)); 
C_55_S_2_L_3_inst : LUT6 generic map(INIT => "1111111100011111011100011011001100000100000001100000000000100001") port map( O =>C_55_S_2_L_3_out, I0 =>  inp_feat(509), I1 =>  inp_feat(334), I2 =>  inp_feat(227), I3 =>  inp_feat(311), I4 =>  inp_feat(476), I5 =>  inp_feat(344)); 
C_55_S_2_L_4_inst : LUT6 generic map(INIT => "1000001100000000101000001001010000000000000000000000000011001000") port map( O =>C_55_S_2_L_4_out, I0 =>  inp_feat(160), I1 =>  inp_feat(178), I2 =>  inp_feat(464), I3 =>  inp_feat(221), I4 =>  inp_feat(74), I5 =>  inp_feat(20)); 
C_55_S_2_L_5_inst : LUT6 generic map(INIT => "0000000000110001000000000000010010101101101101001000000100000010") port map( O =>C_55_S_2_L_5_out, I0 =>  inp_feat(30), I1 =>  inp_feat(96), I2 =>  inp_feat(191), I3 =>  inp_feat(384), I4 =>  inp_feat(281), I5 =>  inp_feat(359)); 
C_55_S_3_L_0_inst : LUT6 generic map(INIT => "0101010000000001110001000000000010000000000000001100010000000000") port map( O =>C_55_S_3_L_0_out, I0 =>  inp_feat(221), I1 =>  inp_feat(272), I2 =>  inp_feat(285), I3 =>  inp_feat(481), I4 =>  inp_feat(255), I5 =>  inp_feat(219)); 
C_55_S_3_L_1_inst : LUT6 generic map(INIT => "1111011101101100001011110000000100000000000000000001011000000000") port map( O =>C_55_S_3_L_1_out, I0 =>  inp_feat(445), I1 =>  inp_feat(446), I2 =>  inp_feat(485), I3 =>  inp_feat(72), I4 =>  inp_feat(401), I5 =>  inp_feat(228)); 
C_55_S_3_L_2_inst : LUT6 generic map(INIT => "0100001001001010010001100001101000000000000000100000001000010111") port map( O =>C_55_S_3_L_2_out, I0 =>  inp_feat(26), I1 =>  inp_feat(257), I2 =>  inp_feat(387), I3 =>  inp_feat(74), I4 =>  inp_feat(432), I5 =>  inp_feat(20)); 
C_55_S_3_L_3_inst : LUT6 generic map(INIT => "1110001011011010011101010000000000000000000000000111000000000000") port map( O =>C_55_S_3_L_3_out, I0 =>  inp_feat(387), I1 =>  inp_feat(231), I2 =>  inp_feat(288), I3 =>  inp_feat(419), I4 =>  inp_feat(432), I5 =>  inp_feat(20)); 
C_55_S_3_L_4_inst : LUT6 generic map(INIT => "0000001010001001000000000011100010101110000011100000000000100000") port map( O =>C_55_S_3_L_4_out, I0 =>  inp_feat(476), I1 =>  inp_feat(133), I2 =>  inp_feat(395), I3 =>  inp_feat(104), I4 =>  inp_feat(40), I5 =>  inp_feat(422)); 
C_55_S_3_L_5_inst : LUT6 generic map(INIT => "0011010011010000010100101101000010101000000000000000000000000000") port map( O =>C_55_S_3_L_5_out, I0 =>  inp_feat(323), I1 =>  inp_feat(387), I2 =>  inp_feat(406), I3 =>  inp_feat(440), I4 =>  inp_feat(306), I5 =>  inp_feat(498)); 
C_55_S_4_L_0_inst : LUT6 generic map(INIT => "1001010101000001110100110000001100000000000001001101001000000000") port map( O =>C_55_S_4_L_0_out, I0 =>  inp_feat(450), I1 =>  inp_feat(49), I2 =>  inp_feat(92), I3 =>  inp_feat(275), I4 =>  inp_feat(160), I5 =>  inp_feat(437)); 
C_55_S_4_L_1_inst : LUT6 generic map(INIT => "0000000000001010000000000000100010101001100010001010000000000000") port map( O =>C_55_S_4_L_1_out, I0 =>  inp_feat(214), I1 =>  inp_feat(160), I2 =>  inp_feat(157), I3 =>  inp_feat(501), I4 =>  inp_feat(197), I5 =>  inp_feat(204)); 
C_55_S_4_L_2_inst : LUT6 generic map(INIT => "0101100110101001010011110000011100000001001001010000000110000001") port map( O =>C_55_S_4_L_2_out, I0 =>  inp_feat(379), I1 =>  inp_feat(312), I2 =>  inp_feat(173), I3 =>  inp_feat(90), I4 =>  inp_feat(98), I5 =>  inp_feat(428)); 
C_55_S_4_L_3_inst : LUT6 generic map(INIT => "1101001000011000000000000000001101010010000000000101000011011111") port map( O =>C_55_S_4_L_3_out, I0 =>  inp_feat(432), I1 =>  inp_feat(263), I2 =>  inp_feat(454), I3 =>  inp_feat(350), I4 =>  inp_feat(397), I5 =>  inp_feat(154)); 
C_55_S_4_L_4_inst : LUT6 generic map(INIT => "0000001100100011011010010001110100010110110110110000100000010000") port map( O =>C_55_S_4_L_4_out, I0 =>  inp_feat(316), I1 =>  inp_feat(253), I2 =>  inp_feat(123), I3 =>  inp_feat(412), I4 =>  inp_feat(461), I5 =>  inp_feat(388)); 
C_55_S_4_L_5_inst : LUT6 generic map(INIT => "1110110111011111001100001011011100010000000000000001011111010111") port map( O =>C_55_S_4_L_5_out, I0 =>  inp_feat(312), I1 =>  inp_feat(432), I2 =>  inp_feat(379), I3 =>  inp_feat(104), I4 =>  inp_feat(316), I5 =>  inp_feat(430)); 
C_55_S_5_L_0_inst : LUT6 generic map(INIT => "0000001000101110001001101010111100000000000010100100100000001111") port map( O =>C_55_S_5_L_0_out, I0 =>  inp_feat(81), I1 =>  inp_feat(425), I2 =>  inp_feat(312), I3 =>  inp_feat(418), I4 =>  inp_feat(387), I5 =>  inp_feat(302)); 
C_55_S_5_L_1_inst : LUT6 generic map(INIT => "1111101100111000000100110001100100010001000000000001000110010001") port map( O =>C_55_S_5_L_1_out, I0 =>  inp_feat(316), I1 =>  inp_feat(432), I2 =>  inp_feat(296), I3 =>  inp_feat(60), I4 =>  inp_feat(98), I5 =>  inp_feat(428)); 
C_55_S_5_L_2_inst : LUT6 generic map(INIT => "0001010110100101100100100000110000000000000000010100000000000000") port map( O =>C_55_S_5_L_2_out, I0 =>  inp_feat(139), I1 =>  inp_feat(238), I2 =>  inp_feat(196), I3 =>  inp_feat(21), I4 =>  inp_feat(493), I5 =>  inp_feat(11)); 
C_55_S_5_L_3_inst : LUT6 generic map(INIT => "0001010001010010101000010000010011101101000011010000000000001000") port map( O =>C_55_S_5_L_3_out, I0 =>  inp_feat(292), I1 =>  inp_feat(97), I2 =>  inp_feat(379), I3 =>  inp_feat(304), I4 =>  inp_feat(22), I5 =>  inp_feat(326)); 
C_55_S_5_L_4_inst : LUT6 generic map(INIT => "0000100001000000110001100100101001110010111100000010100100000000") port map( O =>C_55_S_5_L_4_out, I0 =>  inp_feat(461), I1 =>  inp_feat(126), I2 =>  inp_feat(162), I3 =>  inp_feat(244), I4 =>  inp_feat(16), I5 =>  inp_feat(250)); 
C_55_S_5_L_5_inst : LUT6 generic map(INIT => "1111011010111100010101000111100000000000010001100000100000100100") port map( O =>C_55_S_5_L_5_out, I0 =>  inp_feat(509), I1 =>  inp_feat(510), I2 =>  inp_feat(399), I3 =>  inp_feat(422), I4 =>  inp_feat(440), I5 =>  inp_feat(293)); 
C_56_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000010001011100000001000001110001011101111111") port map( O =>C_56_S_0_L_0_out, I0 =>  inp_feat(151), I1 =>  inp_feat(312), I2 =>  inp_feat(173), I3 =>  inp_feat(221), I4 =>  inp_feat(379), I5 =>  inp_feat(316)); 
C_56_S_0_L_1_inst : LUT6 generic map(INIT => "0000000100010111000100110111111110101001100111111000100100010111") port map( O =>C_56_S_0_L_1_out, I0 =>  inp_feat(312), I1 =>  inp_feat(432), I2 =>  inp_feat(221), I3 =>  inp_feat(173), I4 =>  inp_feat(338), I5 =>  inp_feat(489)); 
C_56_S_0_L_2_inst : LUT6 generic map(INIT => "1111110111100011000010011001000101001100010011010000010100011111") port map( O =>C_56_S_0_L_2_out, I0 =>  inp_feat(257), I1 =>  inp_feat(50), I2 =>  inp_feat(318), I3 =>  inp_feat(81), I4 =>  inp_feat(344), I5 =>  inp_feat(473)); 
C_56_S_0_L_3_inst : LUT6 generic map(INIT => "1011001000100101101000111001111100100010000101110001010101111111") port map( O =>C_56_S_0_L_3_out, I0 =>  inp_feat(221), I1 =>  inp_feat(257), I2 =>  inp_feat(316), I3 =>  inp_feat(418), I4 =>  inp_feat(312), I5 =>  inp_feat(164)); 
C_56_S_0_L_4_inst : LUT6 generic map(INIT => "0100000000101010000000000010101000000000000000100000000000000010") port map( O =>C_56_S_0_L_4_out, I0 =>  inp_feat(227), I1 =>  inp_feat(74), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(256), I5 =>  inp_feat(238)); 
C_56_S_0_L_5_inst : LUT6 generic map(INIT => "1100000101001101000101010101111110000000000000000000000100010111") port map( O =>C_56_S_0_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(432), I2 =>  inp_feat(379), I3 =>  inp_feat(436), I4 =>  inp_feat(282), I5 =>  inp_feat(194)); 
C_56_S_1_L_0_inst : LUT6 generic map(INIT => "0000000100010111000100110111111110101001100111111000100100010111") port map( O =>C_56_S_1_L_0_out, I0 =>  inp_feat(312), I1 =>  inp_feat(432), I2 =>  inp_feat(221), I3 =>  inp_feat(173), I4 =>  inp_feat(338), I5 =>  inp_feat(489)); 
C_56_S_1_L_1_inst : LUT6 generic map(INIT => "1111110111100011000010011001000101001100010011010000010100011111") port map( O =>C_56_S_1_L_1_out, I0 =>  inp_feat(257), I1 =>  inp_feat(50), I2 =>  inp_feat(318), I3 =>  inp_feat(81), I4 =>  inp_feat(344), I5 =>  inp_feat(473)); 
C_56_S_1_L_2_inst : LUT6 generic map(INIT => "1011001000100101101000111001111100100010000101110001010101111111") port map( O =>C_56_S_1_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(257), I2 =>  inp_feat(316), I3 =>  inp_feat(418), I4 =>  inp_feat(312), I5 =>  inp_feat(164)); 
C_56_S_1_L_3_inst : LUT6 generic map(INIT => "0100000000101010000000000010101000000000000000100000000000000010") port map( O =>C_56_S_1_L_3_out, I0 =>  inp_feat(227), I1 =>  inp_feat(74), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(256), I5 =>  inp_feat(238)); 
C_56_S_1_L_4_inst : LUT6 generic map(INIT => "1100000101001101000101010101111110000000000000000000000100010111") port map( O =>C_56_S_1_L_4_out, I0 =>  inp_feat(316), I1 =>  inp_feat(432), I2 =>  inp_feat(379), I3 =>  inp_feat(436), I4 =>  inp_feat(282), I5 =>  inp_feat(194)); 
C_56_S_1_L_5_inst : LUT6 generic map(INIT => "0000011011001010000000101100110000000000000011100000100000001000") port map( O =>C_56_S_1_L_5_out, I0 =>  inp_feat(13), I1 =>  inp_feat(106), I2 =>  inp_feat(404), I3 =>  inp_feat(436), I4 =>  inp_feat(256), I5 =>  inp_feat(238)); 
C_56_S_2_L_0_inst : LUT6 generic map(INIT => "1110100101010100001001110000010010001100010011000100110011001101") port map( O =>C_56_S_2_L_0_out, I0 =>  inp_feat(74), I1 =>  inp_feat(249), I2 =>  inp_feat(257), I3 =>  inp_feat(170), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_56_S_2_L_1_inst : LUT6 generic map(INIT => "0010100000000011001100010001010110110011001001111001111101111111") port map( O =>C_56_S_2_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(257), I2 =>  inp_feat(170), I3 =>  inp_feat(282), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_56_S_2_L_2_inst : LUT6 generic map(INIT => "1010001101010111000100110011111100100000010000010000000000010111") port map( O =>C_56_S_2_L_2_out, I0 =>  inp_feat(372), I1 =>  inp_feat(170), I2 =>  inp_feat(387), I3 =>  inp_feat(316), I4 =>  inp_feat(15), I5 =>  inp_feat(90)); 
C_56_S_2_L_3_inst : LUT6 generic map(INIT => "0111100000000001100100000001000000000001000000000000000000000000") port map( O =>C_56_S_2_L_3_out, I0 =>  inp_feat(376), I1 =>  inp_feat(362), I2 =>  inp_feat(432), I3 =>  inp_feat(303), I4 =>  inp_feat(49), I5 =>  inp_feat(344)); 
C_56_S_2_L_4_inst : LUT6 generic map(INIT => "1111101010100010000000100011101101101110000000110000001000000010") port map( O =>C_56_S_2_L_4_out, I0 =>  inp_feat(194), I1 =>  inp_feat(170), I2 =>  inp_feat(316), I3 =>  inp_feat(282), I4 =>  inp_feat(432), I5 =>  inp_feat(187)); 
C_56_S_2_L_5_inst : LUT6 generic map(INIT => "0000000000000001001101010101011100100011100101110001111101111111") port map( O =>C_56_S_2_L_5_out, I0 =>  inp_feat(387), I1 =>  inp_feat(316), I2 =>  inp_feat(221), I3 =>  inp_feat(253), I4 =>  inp_feat(257), I5 =>  inp_feat(270)); 
C_56_S_3_L_0_inst : LUT6 generic map(INIT => "1101000100010101111110110001011101000101000000111010100100010001") port map( O =>C_56_S_3_L_0_out, I0 =>  inp_feat(221), I1 =>  inp_feat(15), I2 =>  inp_feat(372), I3 =>  inp_feat(391), I4 =>  inp_feat(393), I5 =>  inp_feat(176)); 
C_56_S_3_L_1_inst : LUT6 generic map(INIT => "1010000000000010000010101000101000100000001010110010111010101111") port map( O =>C_56_S_3_L_1_out, I0 =>  inp_feat(450), I1 =>  inp_feat(74), I2 =>  inp_feat(221), I3 =>  inp_feat(316), I4 =>  inp_feat(257), I5 =>  inp_feat(270)); 
C_56_S_3_L_2_inst : LUT6 generic map(INIT => "0000011000100100000011000000110010000100110011010100110011001101") port map( O =>C_56_S_3_L_2_out, I0 =>  inp_feat(312), I1 =>  inp_feat(206), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_3_L_3_inst : LUT6 generic map(INIT => "1100001010000001010000010001001100011111111111110001011101111111") port map( O =>C_56_S_3_L_3_out, I0 =>  inp_feat(257), I1 =>  inp_feat(170), I2 =>  inp_feat(436), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_3_L_4_inst : LUT6 generic map(INIT => "0000001110000001101010110001001110000101011111110011111111111111") port map( O =>C_56_S_3_L_4_out, I0 =>  inp_feat(334), I1 =>  inp_feat(170), I2 =>  inp_feat(436), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_3_L_5_inst : LUT6 generic map(INIT => "1100001010000010100010100010001001000110101010100101101010111010") port map( O =>C_56_S_3_L_5_out, I0 =>  inp_feat(389), I1 =>  inp_feat(170), I2 =>  inp_feat(436), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_4_L_0_inst : LUT6 generic map(INIT => "0100000100000001001000010000001110010011100111110001011101111111") port map( O =>C_56_S_4_L_0_out, I0 =>  inp_feat(248), I1 =>  inp_feat(221), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_4_L_1_inst : LUT6 generic map(INIT => "1011000111000111100101111101111111000001000101010000011100011101") port map( O =>C_56_S_4_L_1_out, I0 =>  inp_feat(316), I1 =>  inp_feat(292), I2 =>  inp_feat(379), I3 =>  inp_feat(257), I4 =>  inp_feat(266), I5 =>  inp_feat(489)); 
C_56_S_4_L_2_inst : LUT6 generic map(INIT => "0010000000000001100111010111011110100011100101110001111101111111") port map( O =>C_56_S_4_L_2_out, I0 =>  inp_feat(387), I1 =>  inp_feat(316), I2 =>  inp_feat(221), I3 =>  inp_feat(253), I4 =>  inp_feat(257), I5 =>  inp_feat(270)); 
C_56_S_4_L_3_inst : LUT6 generic map(INIT => "1110000000011010010000100010101000001000010000100000000001001010") port map( O =>C_56_S_4_L_3_out, I0 =>  inp_feat(121), I1 =>  inp_feat(432), I2 =>  inp_feat(170), I3 =>  inp_feat(312), I4 =>  inp_feat(435), I5 =>  inp_feat(440)); 
C_56_S_4_L_4_inst : LUT6 generic map(INIT => "1100000001001111010001100010111100000000000010100010101010101011") port map( O =>C_56_S_4_L_4_out, I0 =>  inp_feat(480), I1 =>  inp_feat(104), I2 =>  inp_feat(257), I3 =>  inp_feat(316), I4 =>  inp_feat(312), I5 =>  inp_feat(164)); 
C_56_S_4_L_5_inst : LUT6 generic map(INIT => "0011001000010000000110110000000010111010101010000001101000000001") port map( O =>C_56_S_4_L_5_out, I0 =>  inp_feat(26), I1 =>  inp_feat(432), I2 =>  inp_feat(257), I3 =>  inp_feat(249), I4 =>  inp_feat(248), I5 =>  inp_feat(69)); 
C_56_S_5_L_0_inst : LUT6 generic map(INIT => "1100011001000100100001000000110010001100110011010100110011001101") port map( O =>C_56_S_5_L_0_out, I0 =>  inp_feat(312), I1 =>  inp_feat(206), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_5_L_1_inst : LUT6 generic map(INIT => "0000110001000100000011100000110011100100110011010100110011001101") port map( O =>C_56_S_5_L_1_out, I0 =>  inp_feat(312), I1 =>  inp_feat(206), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(270), I5 =>  inp_feat(316)); 
C_56_S_5_L_2_inst : LUT6 generic map(INIT => "0110011010110000001011001010001011111110101110110010000011110010") port map( O =>C_56_S_5_L_2_out, I0 =>  inp_feat(94), I1 =>  inp_feat(121), I2 =>  inp_feat(130), I3 =>  inp_feat(251), I4 =>  inp_feat(182), I5 =>  inp_feat(353)); 
C_56_S_5_L_3_inst : LUT6 generic map(INIT => "1111111111100110101000100010001000000010011001000111001001100010") port map( O =>C_56_S_5_L_3_out, I0 =>  inp_feat(312), I1 =>  inp_feat(353), I2 =>  inp_feat(395), I3 =>  inp_feat(266), I4 =>  inp_feat(188), I5 =>  inp_feat(182)); 
C_56_S_5_L_4_inst : LUT6 generic map(INIT => "0010101100101010001010010000110000101100010011000100110011011101") port map( O =>C_56_S_5_L_4_out, I0 =>  inp_feat(130), I1 =>  inp_feat(510), I2 =>  inp_feat(70), I3 =>  inp_feat(170), I4 =>  inp_feat(418), I5 =>  inp_feat(312)); 
C_56_S_5_L_5_inst : LUT6 generic map(INIT => "1111110100000001100011001000000000010001000000001100000000000000") port map( O =>C_56_S_5_L_5_out, I0 =>  inp_feat(221), I1 =>  inp_feat(248), I2 =>  inp_feat(284), I3 =>  inp_feat(201), I4 =>  inp_feat(394), I5 =>  inp_feat(359)); 
C_57_S_0_L_0_inst : LUT6 generic map(INIT => "1111111111111110111111101110101011111110111010001110000010000000") port map( O =>C_57_S_0_L_0_out, I0 =>  inp_feat(173), I1 =>  inp_feat(312), I2 =>  inp_feat(248), I3 =>  inp_feat(221), I4 =>  inp_feat(379), I5 =>  inp_feat(316)); 
C_57_S_0_L_1_inst : LUT6 generic map(INIT => "1111111100101111111110101111000000011100001111101010101000101000") port map( O =>C_57_S_0_L_1_out, I0 =>  inp_feat(160), I1 =>  inp_feat(71), I2 =>  inp_feat(50), I3 =>  inp_feat(282), I4 =>  inp_feat(464), I5 =>  inp_feat(76)); 
C_57_S_0_L_2_inst : LUT6 generic map(INIT => "1001110111111011011111111111111100011111111111110101011111111111") port map( O =>C_57_S_0_L_2_out, I0 =>  inp_feat(0), I1 =>  inp_feat(29), I2 =>  inp_feat(176), I3 =>  inp_feat(455), I4 =>  inp_feat(292), I5 =>  inp_feat(432)); 
C_57_S_0_L_3_inst : LUT6 generic map(INIT => "0111011111011101111111111111111011111111111111111111111101110111") port map( O =>C_57_S_0_L_3_out, I0 =>  inp_feat(472), I1 =>  inp_feat(306), I2 =>  inp_feat(156), I3 =>  inp_feat(344), I4 =>  inp_feat(487), I5 =>  inp_feat(37)); 
C_57_S_0_L_4_inst : LUT6 generic map(INIT => "1111111011110011111111111111111100101111111111101110111011111111") port map( O =>C_57_S_0_L_4_out, I0 =>  inp_feat(130), I1 =>  inp_feat(205), I2 =>  inp_feat(486), I3 =>  inp_feat(29), I4 =>  inp_feat(480), I5 =>  inp_feat(170)); 
C_57_S_0_L_5_inst : LUT6 generic map(INIT => "0001100110010001101111110011000111111111111111111011111000001011") port map( O =>C_57_S_0_L_5_out, I0 =>  inp_feat(257), I1 =>  inp_feat(445), I2 =>  inp_feat(1), I3 =>  inp_feat(446), I4 =>  inp_feat(282), I5 =>  inp_feat(317)); 
C_57_S_1_L_0_inst : LUT6 generic map(INIT => "1111111100101111111110101111000000011100001111101010101000101000") port map( O =>C_57_S_1_L_0_out, I0 =>  inp_feat(160), I1 =>  inp_feat(71), I2 =>  inp_feat(50), I3 =>  inp_feat(282), I4 =>  inp_feat(464), I5 =>  inp_feat(76)); 
C_57_S_1_L_1_inst : LUT6 generic map(INIT => "1001110111111011011111111111111100011111111111110101011111111111") port map( O =>C_57_S_1_L_1_out, I0 =>  inp_feat(0), I1 =>  inp_feat(29), I2 =>  inp_feat(176), I3 =>  inp_feat(455), I4 =>  inp_feat(292), I5 =>  inp_feat(432)); 
C_57_S_1_L_2_inst : LUT6 generic map(INIT => "0111011111011101111111111111111011111111111111111111111101110111") port map( O =>C_57_S_1_L_2_out, I0 =>  inp_feat(472), I1 =>  inp_feat(306), I2 =>  inp_feat(156), I3 =>  inp_feat(344), I4 =>  inp_feat(487), I5 =>  inp_feat(37)); 
C_57_S_1_L_3_inst : LUT6 generic map(INIT => "1111111011110011111111111111111100101111111111101110111011111111") port map( O =>C_57_S_1_L_3_out, I0 =>  inp_feat(130), I1 =>  inp_feat(205), I2 =>  inp_feat(486), I3 =>  inp_feat(29), I4 =>  inp_feat(480), I5 =>  inp_feat(170)); 
C_57_S_1_L_4_inst : LUT6 generic map(INIT => "0001100110010001101111110011000111111111111111111011111000001011") port map( O =>C_57_S_1_L_4_out, I0 =>  inp_feat(257), I1 =>  inp_feat(445), I2 =>  inp_feat(1), I3 =>  inp_feat(446), I4 =>  inp_feat(282), I5 =>  inp_feat(317)); 
C_57_S_1_L_5_inst : LUT6 generic map(INIT => "1110110111111001111111101111110001111010111110000100001010001000") port map( O =>C_57_S_1_L_5_out, I0 =>  inp_feat(443), I1 =>  inp_feat(448), I2 =>  inp_feat(204), I3 =>  inp_feat(66), I4 =>  inp_feat(301), I5 =>  inp_feat(184)); 
C_57_S_2_L_0_inst : LUT6 generic map(INIT => "1111101011101000111111101100110001011000111010001111100011100000") port map( O =>C_57_S_2_L_0_out, I0 =>  inp_feat(316), I1 =>  inp_feat(387), I2 =>  inp_feat(432), I3 =>  inp_feat(326), I4 =>  inp_feat(50), I5 =>  inp_feat(314)); 
C_57_S_2_L_1_inst : LUT6 generic map(INIT => "0010001010001111111111111010001111111110111011001111111011101000") port map( O =>C_57_S_2_L_1_out, I0 =>  inp_feat(432), I1 =>  inp_feat(289), I2 =>  inp_feat(299), I3 =>  inp_feat(326), I4 =>  inp_feat(50), I5 =>  inp_feat(464)); 
C_57_S_2_L_2_inst : LUT6 generic map(INIT => "1110111111001000111111111101100011101110111000000101110000001000") port map( O =>C_57_S_2_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(74), I2 =>  inp_feat(232), I3 =>  inp_feat(506), I4 =>  inp_feat(91), I5 =>  inp_feat(184)); 
C_57_S_2_L_3_inst : LUT6 generic map(INIT => "0011000011110010101000101110001011110110111111000100101011000100") port map( O =>C_57_S_2_L_3_out, I0 =>  inp_feat(292), I1 =>  inp_feat(272), I2 =>  inp_feat(318), I3 =>  inp_feat(180), I4 =>  inp_feat(506), I5 =>  inp_feat(319)); 
C_57_S_2_L_4_inst : LUT6 generic map(INIT => "1010011110101110101111111101110010100110010000101111001101000000") port map( O =>C_57_S_2_L_4_out, I0 =>  inp_feat(506), I1 =>  inp_feat(493), I2 =>  inp_feat(389), I3 =>  inp_feat(229), I4 =>  inp_feat(479), I5 =>  inp_feat(34)); 
C_57_S_2_L_5_inst : LUT6 generic map(INIT => "1100111011001010000111101011111110001100011001111110010110111111") port map( O =>C_57_S_2_L_5_out, I0 =>  inp_feat(316), I1 =>  inp_feat(387), I2 =>  inp_feat(25), I3 =>  inp_feat(61), I4 =>  inp_feat(91), I5 =>  inp_feat(154)); 
C_57_S_3_L_0_inst : LUT6 generic map(INIT => "1111011110110011111111101110011011111110111011101110111011000010") port map( O =>C_57_S_3_L_0_out, I0 =>  inp_feat(23), I1 =>  inp_feat(401), I2 =>  inp_feat(18), I3 =>  inp_feat(344), I4 =>  inp_feat(487), I5 =>  inp_feat(37)); 
C_57_S_3_L_1_inst : LUT6 generic map(INIT => "0000010111111101111011101111001111111111111111101110111010100010") port map( O =>C_57_S_3_L_1_out, I0 =>  inp_feat(401), I1 =>  inp_feat(1), I2 =>  inp_feat(18), I3 =>  inp_feat(456), I4 =>  inp_feat(487), I5 =>  inp_feat(37)); 
C_57_S_3_L_2_inst : LUT6 generic map(INIT => "1101111111101110111111111111011000101011111010111111111110111010") port map( O =>C_57_S_3_L_2_out, I0 =>  inp_feat(221), I1 =>  inp_feat(325), I2 =>  inp_feat(479), I3 =>  inp_feat(96), I4 =>  inp_feat(249), I5 =>  inp_feat(74)); 
C_57_S_3_L_3_inst : LUT6 generic map(INIT => "1011100101111101101111111111111000101011111001101111111111100111") port map( O =>C_57_S_3_L_3_out, I0 =>  inp_feat(130), I1 =>  inp_feat(111), I2 =>  inp_feat(109), I3 =>  inp_feat(125), I4 =>  inp_feat(11), I5 =>  inp_feat(184)); 
C_57_S_3_L_4_inst : LUT6 generic map(INIT => "0011110101111100111101011111010011111101100110011001000011010000") port map( O =>C_57_S_3_L_4_out, I0 =>  inp_feat(361), I1 =>  inp_feat(387), I2 =>  inp_feat(436), I3 =>  inp_feat(184), I4 =>  inp_feat(257), I5 =>  inp_feat(292)); 
C_57_S_3_L_5_inst : LUT6 generic map(INIT => "1111100011111110101001101111111011000100111110111000100011110010") port map( O =>C_57_S_3_L_5_out, I0 =>  inp_feat(170), I1 =>  inp_feat(387), I2 =>  inp_feat(375), I3 =>  inp_feat(454), I4 =>  inp_feat(257), I5 =>  inp_feat(292)); 
C_57_S_4_L_0_inst : LUT6 generic map(INIT => "1011111111100101111111111010111111111111111111010011100111100010") port map( O =>C_57_S_4_L_0_out, I0 =>  inp_feat(413), I1 =>  inp_feat(174), I2 =>  inp_feat(156), I3 =>  inp_feat(483), I4 =>  inp_feat(417), I5 =>  inp_feat(344)); 
C_57_S_4_L_1_inst : LUT6 generic map(INIT => "0000101000101000111111111100100010101010101010001010111110000000") port map( O =>C_57_S_4_L_1_out, I0 =>  inp_feat(74), I1 =>  inp_feat(316), I2 =>  inp_feat(289), I3 =>  inp_feat(387), I4 =>  inp_feat(84), I5 =>  inp_feat(390)); 
C_57_S_4_L_2_inst : LUT6 generic map(INIT => "0111110111101100111111101011111000111100111011001111111111100000") port map( O =>C_57_S_4_L_2_out, I0 =>  inp_feat(509), I1 =>  inp_feat(210), I2 =>  inp_feat(228), I3 =>  inp_feat(108), I4 =>  inp_feat(389), I5 =>  inp_feat(432)); 
C_57_S_4_L_3_inst : LUT6 generic map(INIT => "1001110011111111111100001110100011011111111110101111111110000000") port map( O =>C_57_S_4_L_3_out, I0 =>  inp_feat(282), I1 =>  inp_feat(108), I2 =>  inp_feat(187), I3 =>  inp_feat(478), I4 =>  inp_feat(184), I5 =>  inp_feat(251)); 
C_57_S_4_L_4_inst : LUT6 generic map(INIT => "0001101111111010111111001111100011101111111101011111111110100000") port map( O =>C_57_S_4_L_4_out, I0 =>  inp_feat(483), I1 =>  inp_feat(476), I2 =>  inp_feat(187), I3 =>  inp_feat(478), I4 =>  inp_feat(184), I5 =>  inp_feat(251)); 
C_57_S_4_L_5_inst : LUT6 generic map(INIT => "1111111111101100111101101110100011111111100010000101101010000000") port map( O =>C_57_S_4_L_5_out, I0 =>  inp_feat(379), I1 =>  inp_feat(170), I2 =>  inp_feat(432), I3 =>  inp_feat(316), I4 =>  inp_feat(338), I5 =>  inp_feat(326)); 
C_57_S_5_L_0_inst : LUT6 generic map(INIT => "1101001100101111111111111100011011011111111010111111111111111111") port map( O =>C_57_S_5_L_0_out, I0 =>  inp_feat(200), I1 =>  inp_feat(378), I2 =>  inp_feat(263), I3 =>  inp_feat(72), I4 =>  inp_feat(322), I5 =>  inp_feat(377)); 
C_57_S_5_L_1_inst : LUT6 generic map(INIT => "1011101011111101111111111111100011101000111010001010000010001000") port map( O =>C_57_S_5_L_1_out, I0 =>  inp_feat(143), I1 =>  inp_feat(178), I2 =>  inp_feat(0), I3 =>  inp_feat(263), I4 =>  inp_feat(377), I5 =>  inp_feat(390)); 
C_57_S_5_L_2_inst : LUT6 generic map(INIT => "0000011011111010001011110111110011111111011110110111111111111111") port map( O =>C_57_S_5_L_2_out, I0 =>  inp_feat(45), I1 =>  inp_feat(397), I2 =>  inp_feat(448), I3 =>  inp_feat(65), I4 =>  inp_feat(322), I5 =>  inp_feat(377)); 
C_57_S_5_L_3_inst : LUT6 generic map(INIT => "1111011011110111100011101111111011111111111111100110100011111101") port map( O =>C_57_S_5_L_3_out, I0 =>  inp_feat(316), I1 =>  inp_feat(170), I2 =>  inp_feat(187), I3 =>  inp_feat(92), I4 =>  inp_feat(74), I5 =>  inp_feat(38)); 
C_57_S_5_L_4_inst : LUT6 generic map(INIT => "0010111000111111110111111111111111111000101010101010100010001100") port map( O =>C_57_S_5_L_4_out, I0 =>  inp_feat(106), I1 =>  inp_feat(21), I2 =>  inp_feat(105), I3 =>  inp_feat(180), I4 =>  inp_feat(319), I5 =>  inp_feat(390)); 
C_57_S_5_L_5_inst : LUT6 generic map(INIT => "1100110111100011111111001010110011111100111111011111010001111100") port map( O =>C_57_S_5_L_5_out, I0 =>  inp_feat(89), I1 =>  inp_feat(312), I2 =>  inp_feat(93), I3 =>  inp_feat(407), I4 =>  inp_feat(238), I5 =>  inp_feat(94)); 
C_58_S_0_L_0_inst : LUT6 generic map(INIT => "0000000000000001000000000001001100000001000101110001111101111111") port map( O =>C_58_S_0_L_0_out, I0 =>  inp_feat(312), I1 =>  inp_feat(170), I2 =>  inp_feat(248), I3 =>  inp_feat(221), I4 =>  inp_feat(379), I5 =>  inp_feat(316)); 
C_58_S_0_L_1_inst : LUT6 generic map(INIT => "0001000000001111001101011001111100110011001101111111011111111111") port map( O =>C_58_S_0_L_1_out, I0 =>  inp_feat(253), I1 =>  inp_feat(334), I2 =>  inp_feat(432), I3 =>  inp_feat(257), I4 =>  inp_feat(130), I5 =>  inp_feat(282)); 
C_58_S_0_L_2_inst : LUT6 generic map(INIT => "0111011111100001111000110111010100000000000100010001000001110001") port map( O =>C_58_S_0_L_2_out, I0 =>  inp_feat(316), I1 =>  inp_feat(379), I2 =>  inp_feat(82), I3 =>  inp_feat(170), I4 =>  inp_feat(372), I5 =>  inp_feat(494)); 
C_58_S_0_L_3_inst : LUT6 generic map(INIT => "0011011100011111111001111001011100000001000101010000000100110111") port map( O =>C_58_S_0_L_3_out, I0 =>  inp_feat(387), I1 =>  inp_feat(173), I2 =>  inp_feat(418), I3 =>  inp_feat(221), I4 =>  inp_feat(412), I5 =>  inp_feat(494)); 
C_58_S_0_L_4_inst : LUT6 generic map(INIT => "1111001111011111000000010001010100000000000000000000000000000000") port map( O =>C_58_S_0_L_4_out, I0 =>  inp_feat(312), I1 =>  inp_feat(289), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(494), I5 =>  inp_feat(33)); 
C_58_S_0_L_5_inst : LUT6 generic map(INIT => "0011010100110001001000010000101000111001000100001000001010001010") port map( O =>C_58_S_0_L_5_out, I0 =>  inp_feat(432), I1 =>  inp_feat(338), I2 =>  inp_feat(258), I3 =>  inp_feat(97), I4 =>  inp_feat(288), I5 =>  inp_feat(117)); 
C_58_S_1_L_0_inst : LUT6 generic map(INIT => "0001000000001111001101011001111100110011001101111111011111111111") port map( O =>C_58_S_1_L_0_out, I0 =>  inp_feat(253), I1 =>  inp_feat(334), I2 =>  inp_feat(432), I3 =>  inp_feat(257), I4 =>  inp_feat(130), I5 =>  inp_feat(282)); 
C_58_S_1_L_1_inst : LUT6 generic map(INIT => "0111011111100001111000110111010100000000000100010001000001110001") port map( O =>C_58_S_1_L_1_out, I0 =>  inp_feat(316), I1 =>  inp_feat(379), I2 =>  inp_feat(82), I3 =>  inp_feat(170), I4 =>  inp_feat(372), I5 =>  inp_feat(494)); 
C_58_S_1_L_2_inst : LUT6 generic map(INIT => "0011011100011111111001111001011100000001000101010000000100110111") port map( O =>C_58_S_1_L_2_out, I0 =>  inp_feat(387), I1 =>  inp_feat(173), I2 =>  inp_feat(418), I3 =>  inp_feat(221), I4 =>  inp_feat(412), I5 =>  inp_feat(494)); 
C_58_S_1_L_3_inst : LUT6 generic map(INIT => "1111001111011111000000010001010100000000000000000000000000000000") port map( O =>C_58_S_1_L_3_out, I0 =>  inp_feat(312), I1 =>  inp_feat(289), I2 =>  inp_feat(170), I3 =>  inp_feat(372), I4 =>  inp_feat(494), I5 =>  inp_feat(33)); 
C_58_S_1_L_4_inst : LUT6 generic map(INIT => "0011010100110001001000010000101000111001000100001000001010001010") port map( O =>C_58_S_1_L_4_out, I0 =>  inp_feat(432), I1 =>  inp_feat(338), I2 =>  inp_feat(258), I3 =>  inp_feat(97), I4 =>  inp_feat(288), I5 =>  inp_feat(117)); 
C_58_S_1_L_5_inst : LUT6 generic map(INIT => "1000110101000101000000000010000010101110011111110000100000000110") port map( O =>C_58_S_1_L_5_out, I0 =>  inp_feat(432), I1 =>  inp_feat(307), I2 =>  inp_feat(163), I3 =>  inp_feat(46), I4 =>  inp_feat(437), I5 =>  inp_feat(127)); 
C_58_S_2_L_0_inst : LUT6 generic map(INIT => "0001010100010111010101111111111100000000000101110000000000111111") port map( O =>C_58_S_2_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(418), I2 =>  inp_feat(173), I3 =>  inp_feat(312), I4 =>  inp_feat(130), I5 =>  inp_feat(494)); 
C_58_S_2_L_1_inst : LUT6 generic map(INIT => "1001011010110001110111001111000100000000000000000000000001110000") port map( O =>C_58_S_2_L_1_out, I0 =>  inp_feat(221), I1 =>  inp_feat(257), I2 =>  inp_feat(175), I3 =>  inp_feat(312), I4 =>  inp_feat(248), I5 =>  inp_feat(494)); 
C_58_S_2_L_2_inst : LUT6 generic map(INIT => "0010001100010011111010100000000000000000000000000000001000000000") port map( O =>C_58_S_2_L_2_out, I0 =>  inp_feat(249), I1 =>  inp_feat(151), I2 =>  inp_feat(282), I3 =>  inp_feat(344), I4 =>  inp_feat(368), I5 =>  inp_feat(33)); 
C_58_S_2_L_3_inst : LUT6 generic map(INIT => "0100000111000000101100010000000000000000000000000000000000000000") port map( O =>C_58_S_2_L_3_out, I0 =>  inp_feat(289), I1 =>  inp_feat(99), I2 =>  inp_feat(313), I3 =>  inp_feat(283), I4 =>  inp_feat(116), I5 =>  inp_feat(33)); 
C_58_S_2_L_4_inst : LUT6 generic map(INIT => "0110010110100001001101100000100010011101001101110000010000000000") port map( O =>C_58_S_2_L_4_out, I0 =>  inp_feat(366), I1 =>  inp_feat(445), I2 =>  inp_feat(379), I3 =>  inp_feat(406), I4 =>  inp_feat(305), I5 =>  inp_feat(372)); 
C_58_S_2_L_5_inst : LUT6 generic map(INIT => "1111100100011000101100010000000000000000000000000001111100000010") port map( O =>C_58_S_2_L_5_out, I0 =>  inp_feat(187), I1 =>  inp_feat(163), I2 =>  inp_feat(105), I3 =>  inp_feat(179), I4 =>  inp_feat(123), I5 =>  inp_feat(244)); 
C_58_S_3_L_0_inst : LUT6 generic map(INIT => "0001000001110000101100011111001100000000000000000000000011110010") port map( O =>C_58_S_3_L_0_out, I0 =>  inp_feat(442), I1 =>  inp_feat(104), I2 =>  inp_feat(201), I3 =>  inp_feat(312), I4 =>  inp_feat(173), I5 =>  inp_feat(494)); 
C_58_S_3_L_1_inst : LUT6 generic map(INIT => "0000011110110100100111010011111100000001000000110000001100011011") port map( O =>C_58_S_3_L_1_out, I0 =>  inp_feat(151), I1 =>  inp_feat(316), I2 =>  inp_feat(379), I3 =>  inp_feat(170), I4 =>  inp_feat(372), I5 =>  inp_feat(494)); 
C_58_S_3_L_2_inst : LUT6 generic map(INIT => "1100000001100000101000011011001000000000000000000000000010100010") port map( O =>C_58_S_3_L_2_out, I0 =>  inp_feat(114), I1 =>  inp_feat(104), I2 =>  inp_feat(201), I3 =>  inp_feat(312), I4 =>  inp_feat(173), I5 =>  inp_feat(494)); 
C_58_S_3_L_3_inst : LUT6 generic map(INIT => "0010100100100101111000100000000000000000000000000000000000000000") port map( O =>C_58_S_3_L_3_out, I0 =>  inp_feat(304), I1 =>  inp_feat(115), I2 =>  inp_feat(500), I3 =>  inp_feat(49), I4 =>  inp_feat(474), I5 =>  inp_feat(33)); 
C_58_S_3_L_4_inst : LUT6 generic map(INIT => "1111010100011001000111010001101100110010000000000000110000000000") port map( O =>C_58_S_3_L_4_out, I0 =>  inp_feat(74), I1 =>  inp_feat(356), I2 =>  inp_feat(449), I3 =>  inp_feat(453), I4 =>  inp_feat(460), I5 =>  inp_feat(89)); 
C_58_S_3_L_5_inst : LUT6 generic map(INIT => "0000000100000011000000100000010110110100000000000000000000000000") port map( O =>C_58_S_3_L_5_out, I0 =>  inp_feat(165), I1 =>  inp_feat(412), I2 =>  inp_feat(99), I3 =>  inp_feat(124), I4 =>  inp_feat(419), I5 =>  inp_feat(34)); 
C_58_S_4_L_0_inst : LUT6 generic map(INIT => "1111011100011111101001010010101100000001000000110000000100001101") port map( O =>C_58_S_4_L_0_out, I0 =>  inp_feat(372), I1 =>  inp_feat(418), I2 =>  inp_feat(387), I3 =>  inp_feat(326), I4 =>  inp_feat(255), I5 =>  inp_feat(499)); 
C_58_S_4_L_1_inst : LUT6 generic map(INIT => "0011110010000010100010101111111000000000000000000000000011000010") port map( O =>C_58_S_4_L_1_out, I0 =>  inp_feat(322), I1 =>  inp_feat(190), I2 =>  inp_feat(135), I3 =>  inp_feat(325), I4 =>  inp_feat(133), I5 =>  inp_feat(453)); 
C_58_S_4_L_2_inst : LUT6 generic map(INIT => "0000000000001110011000000000000010101110000011000000000000000100") port map( O =>C_58_S_4_L_2_out, I0 =>  inp_feat(407), I1 =>  inp_feat(300), I2 =>  inp_feat(338), I3 =>  inp_feat(448), I4 =>  inp_feat(153), I5 =>  inp_feat(379)); 
C_58_S_4_L_3_inst : LUT6 generic map(INIT => "1000111110001101110011110000011100000100000000000000000000000000") port map( O =>C_58_S_4_L_3_out, I0 =>  inp_feat(147), I1 =>  inp_feat(489), I2 =>  inp_feat(282), I3 =>  inp_feat(448), I4 =>  inp_feat(84), I5 =>  inp_feat(33)); 
C_58_S_4_L_4_inst : LUT6 generic map(INIT => "0011011111010010000000001010000111111011101000001001000010100000") port map( O =>C_58_S_4_L_4_out, I0 =>  inp_feat(420), I1 =>  inp_feat(160), I2 =>  inp_feat(27), I3 =>  inp_feat(270), I4 =>  inp_feat(384), I5 =>  inp_feat(133)); 
C_58_S_4_L_5_inst : LUT6 generic map(INIT => "0011011100000011100000010010010110011111100000100001110000000000") port map( O =>C_58_S_4_L_5_out, I0 =>  inp_feat(379), I1 =>  inp_feat(115), I2 =>  inp_feat(151), I3 =>  inp_feat(246), I4 =>  inp_feat(448), I5 =>  inp_feat(84)); 
C_58_S_5_L_0_inst : LUT6 generic map(INIT => "1000000000010011000000000000000010110011101100110101000010000011") port map( O =>C_58_S_5_L_0_out, I0 =>  inp_feat(456), I1 =>  inp_feat(108), I2 =>  inp_feat(344), I3 =>  inp_feat(390), I4 =>  inp_feat(437), I5 =>  inp_feat(127)); 
C_58_S_5_L_1_inst : LUT6 generic map(INIT => "0000010100000001000001001000000011101111001011100000000000000010") port map( O =>C_58_S_5_L_1_out, I0 =>  inp_feat(323), I1 =>  inp_feat(385), I2 =>  inp_feat(16), I3 =>  inp_feat(105), I4 =>  inp_feat(124), I5 =>  inp_feat(334)); 
C_58_S_5_L_2_inst : LUT6 generic map(INIT => "0001101010001100001000000000110010001101110011000000000000001110") port map( O =>C_58_S_5_L_2_out, I0 =>  inp_feat(322), I1 =>  inp_feat(195), I2 =>  inp_feat(257), I3 =>  inp_feat(292), I4 =>  inp_feat(507), I5 =>  inp_feat(416)); 
C_58_S_5_L_3_inst : LUT6 generic map(INIT => "0011000011110000000000101000000110010010111100001111111100100100") port map( O =>C_58_S_5_L_3_out, I0 =>  inp_feat(1), I1 =>  inp_feat(331), I2 =>  inp_feat(339), I3 =>  inp_feat(412), I4 =>  inp_feat(226), I5 =>  inp_feat(233)); 
C_58_S_5_L_4_inst : LUT6 generic map(INIT => "1101110100011100100011000000010000100001000001000000010101000000") port map( O =>C_58_S_5_L_4_out, I0 =>  inp_feat(76), I1 =>  inp_feat(299), I2 =>  inp_feat(391), I3 =>  inp_feat(384), I4 =>  inp_feat(474), I5 =>  inp_feat(272)); 
C_58_S_5_L_5_inst : LUT6 generic map(INIT => "0001000010011000000000001100000011110000101011000001000000000000") port map( O =>C_58_S_5_L_5_out, I0 =>  inp_feat(202), I1 =>  inp_feat(48), I2 =>  inp_feat(373), I3 =>  inp_feat(406), I4 =>  inp_feat(305), I5 =>  inp_feat(372)); 
C_59_S_0_L_0_inst : LUT6 generic map(INIT => "1111111011111110111111101110110011111010111010001110000010000000") port map( O =>C_59_S_0_L_0_out, I0 =>  inp_feat(312), I1 =>  inp_feat(170), I2 =>  inp_feat(248), I3 =>  inp_feat(221), I4 =>  inp_feat(379), I5 =>  inp_feat(316)); 
C_59_S_0_L_1_inst : LUT6 generic map(INIT => "0000010000001000111111101000100011111111111010001111010111111111") port map( O =>C_59_S_0_L_1_out, I0 =>  inp_feat(292), I1 =>  inp_feat(387), I2 =>  inp_feat(391), I3 =>  inp_feat(372), I4 =>  inp_feat(10), I5 =>  inp_feat(169)); 
C_59_S_0_L_2_inst : LUT6 generic map(INIT => "1111111111111110100110101110000000111100110110101100100000000000") port map( O =>C_59_S_0_L_2_out, I0 =>  inp_feat(282), I1 =>  inp_feat(391), I2 =>  inp_feat(418), I3 =>  inp_feat(432), I4 =>  inp_feat(387), I5 =>  inp_feat(316)); 
C_59_S_0_L_3_inst : LUT6 generic map(INIT => "1111111001011110111100101110101111111111010011000010001011110001") port map( O =>C_59_S_0_L_3_out, I0 =>  inp_feat(37), I1 =>  inp_feat(104), I2 =>  inp_feat(510), I3 =>  inp_feat(312), I4 =>  inp_feat(91), I5 =>  inp_feat(250)); 
C_59_S_0_L_4_inst : LUT6 generic map(INIT => "1110101111111010000011100001001001101110110110001111110010010000") port map( O =>C_59_S_0_L_4_out, I0 =>  inp_feat(189), I1 =>  inp_feat(8), I2 =>  inp_feat(159), I3 =>  inp_feat(348), I4 =>  inp_feat(11), I5 =>  inp_feat(363)); 
C_59_S_0_L_5_inst : LUT6 generic map(INIT => "1010101110100110011100111111000001101110011010000011001111100000") port map( O =>C_59_S_0_L_5_out, I0 =>  inp_feat(231), I1 =>  inp_feat(454), I2 =>  inp_feat(470), I3 =>  inp_feat(453), I4 =>  inp_feat(263), I5 =>  inp_feat(76)); 
C_59_S_1_L_0_inst : LUT6 generic map(INIT => "0000010000001000111111101000100011111111111010001111010111111111") port map( O =>C_59_S_1_L_0_out, I0 =>  inp_feat(292), I1 =>  inp_feat(387), I2 =>  inp_feat(391), I3 =>  inp_feat(372), I4 =>  inp_feat(10), I5 =>  inp_feat(169)); 
C_59_S_1_L_1_inst : LUT6 generic map(INIT => "1111111111111110100110101110000000111100110110101100100000000000") port map( O =>C_59_S_1_L_1_out, I0 =>  inp_feat(282), I1 =>  inp_feat(391), I2 =>  inp_feat(418), I3 =>  inp_feat(432), I4 =>  inp_feat(387), I5 =>  inp_feat(316)); 
C_59_S_1_L_2_inst : LUT6 generic map(INIT => "1111111001011110111100101110101111111111010011000010001011110001") port map( O =>C_59_S_1_L_2_out, I0 =>  inp_feat(37), I1 =>  inp_feat(104), I2 =>  inp_feat(510), I3 =>  inp_feat(312), I4 =>  inp_feat(91), I5 =>  inp_feat(250)); 
C_59_S_1_L_3_inst : LUT6 generic map(INIT => "1110101111111010000011100001001001101110110110001111110010010000") port map( O =>C_59_S_1_L_3_out, I0 =>  inp_feat(189), I1 =>  inp_feat(8), I2 =>  inp_feat(159), I3 =>  inp_feat(348), I4 =>  inp_feat(11), I5 =>  inp_feat(363)); 
C_59_S_1_L_4_inst : LUT6 generic map(INIT => "1010101110100110011100111111000001101110011010000011001111100000") port map( O =>C_59_S_1_L_4_out, I0 =>  inp_feat(231), I1 =>  inp_feat(454), I2 =>  inp_feat(470), I3 =>  inp_feat(453), I4 =>  inp_feat(263), I5 =>  inp_feat(76)); 
C_59_S_1_L_5_inst : LUT6 generic map(INIT => "1101111101100111110011110011110011111111101100100001001100100010") port map( O =>C_59_S_1_L_5_out, I0 =>  inp_feat(292), I1 =>  inp_feat(328), I2 =>  inp_feat(374), I3 =>  inp_feat(379), I4 =>  inp_feat(257), I5 =>  inp_feat(432)); 
C_59_S_2_L_0_inst : LUT6 generic map(INIT => "1100001111111010111011101100100000010010011111011111001111111111") port map( O =>C_59_S_2_L_0_out, I0 =>  inp_feat(391), I1 =>  inp_feat(350), I2 =>  inp_feat(387), I3 =>  inp_feat(201), I4 =>  inp_feat(169), I5 =>  inp_feat(379)); 
C_59_S_2_L_1_inst : LUT6 generic map(INIT => "1100110011100110101000001010010001101000111010000010100000101000") port map( O =>C_59_S_2_L_1_out, I0 =>  inp_feat(312), I1 =>  inp_feat(282), I2 =>  inp_feat(74), I3 =>  inp_feat(212), I4 =>  inp_feat(368), I5 =>  inp_feat(463)); 
C_59_S_2_L_2_inst : LUT6 generic map(INIT => "1000101010011000111111000000100001010011111100100111111111001000") port map( O =>C_59_S_2_L_2_out, I0 =>  inp_feat(289), I1 =>  inp_feat(470), I2 =>  inp_feat(432), I3 =>  inp_feat(429), I4 =>  inp_feat(106), I5 =>  inp_feat(300)); 
C_59_S_2_L_3_inst : LUT6 generic map(INIT => "1010000111101011011111101111110010100010000000001111111111011111") port map( O =>C_59_S_2_L_3_out, I0 =>  inp_feat(379), I1 =>  inp_feat(267), I2 =>  inp_feat(63), I3 =>  inp_feat(254), I4 =>  inp_feat(142), I5 =>  inp_feat(224)); 
C_59_S_2_L_4_inst : LUT6 generic map(INIT => "1110110111110001001010111111111000101010110101011111111010111001") port map( O =>C_59_S_2_L_4_out, I0 =>  inp_feat(366), I1 =>  inp_feat(182), I2 =>  inp_feat(472), I3 =>  inp_feat(279), I4 =>  inp_feat(282), I5 =>  inp_feat(244)); 
C_59_S_2_L_5_inst : LUT6 generic map(INIT => "0100000101000110001001011000000011111110110101001110100010000000") port map( O =>C_59_S_2_L_5_out, I0 =>  inp_feat(104), I1 =>  inp_feat(316), I2 =>  inp_feat(418), I3 =>  inp_feat(387), I4 =>  inp_feat(432), I5 =>  inp_feat(282)); 
C_59_S_3_L_0_inst : LUT6 generic map(INIT => "0010100100101001001011101111011111111110111111001100000001110000") port map( O =>C_59_S_3_L_0_out, I0 =>  inp_feat(446), I1 =>  inp_feat(199), I2 =>  inp_feat(108), I3 =>  inp_feat(107), I4 =>  inp_feat(486), I5 =>  inp_feat(20)); 
C_59_S_3_L_1_inst : LUT6 generic map(INIT => "1010011110011110100001100000110111011110111111011100110001000100") port map( O =>C_59_S_3_L_1_out, I0 =>  inp_feat(248), I1 =>  inp_feat(316), I2 =>  inp_feat(374), I3 =>  inp_feat(287), I4 =>  inp_feat(119), I5 =>  inp_feat(304)); 
C_59_S_3_L_2_inst : LUT6 generic map(INIT => "1001101110001001110111010000110011011000110110011010111000001100") port map( O =>C_59_S_3_L_2_out, I0 =>  inp_feat(152), I1 =>  inp_feat(289), I2 =>  inp_feat(287), I3 =>  inp_feat(387), I4 =>  inp_feat(183), I5 =>  inp_feat(304)); 
C_59_S_3_L_3_inst : LUT6 generic map(INIT => "1110110101010111100110000101111101101000001011101010010111110101") port map( O =>C_59_S_3_L_3_out, I0 =>  inp_feat(189), I1 =>  inp_feat(110), I2 =>  inp_feat(176), I3 =>  inp_feat(392), I4 =>  inp_feat(398), I5 =>  inp_feat(106)); 
C_59_S_3_L_4_inst : LUT6 generic map(INIT => "0010000011010001000010111011011111101001101010101000101010000010") port map( O =>C_59_S_3_L_4_out, I0 =>  inp_feat(312), I1 =>  inp_feat(221), I2 =>  inp_feat(91), I3 =>  inp_feat(101), I4 =>  inp_feat(102), I5 =>  inp_feat(266)); 
C_59_S_3_L_5_inst : LUT6 generic map(INIT => "1110111001111100000011100000110111011110111011101100110000000100") port map( O =>C_59_S_3_L_5_out, I0 =>  inp_feat(282), I1 =>  inp_feat(316), I2 =>  inp_feat(374), I3 =>  inp_feat(287), I4 =>  inp_feat(119), I5 =>  inp_feat(304)); 
C_59_S_4_L_0_inst : LUT6 generic map(INIT => "1101110101011100110111011111110111101100101000000000000000101100") port map( O =>C_59_S_4_L_0_out, I0 =>  inp_feat(127), I1 =>  inp_feat(372), I2 =>  inp_feat(253), I3 =>  inp_feat(12), I4 =>  inp_feat(190), I5 =>  inp_feat(88)); 
C_59_S_4_L_1_inst : LUT6 generic map(INIT => "1111001010110011100110011111101000111000111110111111101011111011") port map( O =>C_59_S_4_L_1_out, I0 =>  inp_feat(130), I1 =>  inp_feat(158), I2 =>  inp_feat(368), I3 =>  inp_feat(183), I4 =>  inp_feat(261), I5 =>  inp_feat(47)); 
C_59_S_4_L_2_inst : LUT6 generic map(INIT => "0001001111110111000110111101001111111101111110111101111110101100") port map( O =>C_59_S_4_L_2_out, I0 =>  inp_feat(13), I1 =>  inp_feat(508), I2 =>  inp_feat(491), I3 =>  inp_feat(105), I4 =>  inp_feat(79), I5 =>  inp_feat(81)); 
C_59_S_4_L_3_inst : LUT6 generic map(INIT => "1010000111100111010101001111000000100110110100000110110011100000") port map( O =>C_59_S_4_L_3_out, I0 =>  inp_feat(437), I1 =>  inp_feat(231), I2 =>  inp_feat(123), I3 =>  inp_feat(384), I4 =>  inp_feat(205), I5 =>  inp_feat(474)); 
C_59_S_4_L_4_inst : LUT6 generic map(INIT => "1110101010111010010111111011000110011011001111000100110011001000") port map( O =>C_59_S_4_L_4_out, I0 =>  inp_feat(249), I1 =>  inp_feat(173), I2 =>  inp_feat(108), I3 =>  inp_feat(415), I4 =>  inp_feat(387), I5 =>  inp_feat(432)); 
C_59_S_4_L_5_inst : LUT6 generic map(INIT => "1100111001011101110111110101111101101100010011001111011001100100") port map( O =>C_59_S_4_L_5_out, I0 =>  inp_feat(22), I1 =>  inp_feat(464), I2 =>  inp_feat(426), I3 =>  inp_feat(277), I4 =>  inp_feat(124), I5 =>  inp_feat(486)); 
C_59_S_5_L_0_inst : LUT6 generic map(INIT => "0001111111111101101011100111111011011110111100100000100011000100") port map( O =>C_59_S_5_L_0_out, I0 =>  inp_feat(387), I1 =>  inp_feat(314), I2 =>  inp_feat(421), I3 =>  inp_feat(204), I4 =>  inp_feat(432), I5 =>  inp_feat(282)); 
C_59_S_5_L_1_inst : LUT6 generic map(INIT => "1111101011000011111100110100110000001010010011101111111111111000") port map( O =>C_59_S_5_L_1_out, I0 =>  inp_feat(472), I1 =>  inp_feat(242), I2 =>  inp_feat(465), I3 =>  inp_feat(78), I4 =>  inp_feat(19), I5 =>  inp_feat(72)); 
C_59_S_5_L_2_inst : LUT6 generic map(INIT => "0010000000101101011110100110101010111111111000101111101011101001") port map( O =>C_59_S_5_L_2_out, I0 =>  inp_feat(508), I1 =>  inp_feat(108), I2 =>  inp_feat(486), I3 =>  inp_feat(107), I4 =>  inp_feat(475), I5 =>  inp_feat(39)); 
C_59_S_5_L_3_inst : LUT6 generic map(INIT => "1000101101001101101001111111110011011011001001101111111111111101") port map( O =>C_59_S_5_L_3_out, I0 =>  inp_feat(347), I1 =>  inp_feat(391), I2 =>  inp_feat(392), I3 =>  inp_feat(313), I4 =>  inp_feat(227), I5 =>  inp_feat(371)); 
C_59_S_5_L_4_inst : LUT6 generic map(INIT => "0111000111011010110100100010111111111111111111111111111000011111") port map( O =>C_59_S_5_L_4_out, I0 =>  inp_feat(281), I1 =>  inp_feat(284), I2 =>  inp_feat(258), I3 =>  inp_feat(428), I4 =>  inp_feat(201), I5 =>  inp_feat(220)); 
C_59_S_5_L_5_inst : LUT6 generic map(INIT => "1110110111101010101010000100100001001100001010001111101010100000") port map( O =>C_59_S_5_L_5_out, I0 =>  inp_feat(270), I1 =>  inp_feat(436), I2 =>  inp_feat(212), I3 =>  inp_feat(485), I4 =>  inp_feat(61), I5 =>  inp_feat(254)); 

C_0_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_0_S_0_out, I0 =>  C_0_S_0_L_0_out, I1 =>  C_0_S_0_L_1_out, I2 =>  C_0_S_0_L_2_out, I3 =>  C_0_S_0_L_3_out, I4 =>  C_0_S_0_L_4_out, I5 =>  C_0_S_0_L_5_out); 
C_0_S_1_inst : LUT6 generic map(INIT => "1110101011101010111010101010100011101010101010001010100010101000") port map( O =>C_0_S_1_out, I0 =>  C_0_S_1_L_0_out, I1 =>  C_0_S_1_L_1_out, I2 =>  C_0_S_1_L_2_out, I3 =>  C_0_S_1_L_3_out, I4 =>  C_0_S_1_L_4_out, I5 =>  C_0_S_1_L_5_out); 
C_0_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010101010100011101010101010001110100010000000") port map( O =>C_0_S_2_out, I0 =>  C_0_S_2_L_0_out, I1 =>  C_0_S_2_L_1_out, I2 =>  C_0_S_2_L_2_out, I3 =>  C_0_S_2_L_3_out, I4 =>  C_0_S_2_L_4_out, I5 =>  C_0_S_2_L_5_out); 
C_0_S_3_inst : LUT6 generic map(INIT => "1111111011111110111111001110100011101000110000001000000010000000") port map( O =>C_0_S_3_out, I0 =>  C_0_S_3_L_0_out, I1 =>  C_0_S_3_L_1_out, I2 =>  C_0_S_3_L_2_out, I3 =>  C_0_S_3_L_3_out, I4 =>  C_0_S_3_L_4_out, I5 =>  C_0_S_3_L_5_out); 
C_0_S_4_inst : LUT6 generic map(INIT => "1111111111111010111111101010000011111010100000001010000000000000") port map( O =>C_0_S_4_out, I0 =>  C_0_S_4_L_0_out, I1 =>  C_0_S_4_L_1_out, I2 =>  C_0_S_4_L_2_out, I3 =>  C_0_S_4_L_3_out, I4 =>  C_0_S_4_L_4_out, I5 =>  C_0_S_4_L_5_out); 
C_0_S_5_inst : LUT6 generic map(INIT => "1111111011111000111110101110000011111000101000001110000010000000") port map( O =>C_0_S_5_out, I0 =>  C_0_S_5_L_0_out, I1 =>  C_0_S_5_L_1_out, I2 =>  C_0_S_5_L_2_out, I3 =>  C_0_S_5_L_3_out, I4 =>  C_0_S_5_L_4_out, I5 =>  C_0_S_5_L_5_out); 

C_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_0_out, I0 =>  C_0_S_0_out, I1 =>  C_0_S_1_out, I2 =>  C_0_S_2_out, I3 =>  C_0_S_3_out, I4 =>  C_0_S_4_out, I5 =>  C_0_S_5_out); 

 
C_1_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_1_S_0_out, I0 =>  C_1_S_0_L_0_out, I1 =>  C_1_S_0_L_1_out, I2 =>  C_1_S_0_L_2_out, I3 =>  C_1_S_0_L_3_out, I4 =>  C_1_S_0_L_4_out, I5 =>  C_1_S_0_L_5_out); 
C_1_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_1_S_1_out, I0 =>  C_1_S_1_L_0_out, I1 =>  C_1_S_1_L_1_out, I2 =>  C_1_S_1_L_2_out, I3 =>  C_1_S_1_L_3_out, I4 =>  C_1_S_1_L_4_out, I5 =>  C_1_S_1_L_5_out); 
C_1_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_1_S_2_out, I0 =>  C_1_S_2_L_0_out, I1 =>  C_1_S_2_L_1_out, I2 =>  C_1_S_2_L_2_out, I3 =>  C_1_S_2_L_3_out, I4 =>  C_1_S_2_L_4_out, I5 =>  C_1_S_2_L_5_out); 
C_1_S_3_inst : LUT6 generic map(INIT => "1111111111111100111111001100000011111100110000001100000000000000") port map( O =>C_1_S_3_out, I0 =>  C_1_S_3_L_0_out, I1 =>  C_1_S_3_L_1_out, I2 =>  C_1_S_3_L_2_out, I3 =>  C_1_S_3_L_3_out, I4 =>  C_1_S_3_L_4_out, I5 =>  C_1_S_3_L_5_out); 
C_1_S_4_inst : LUT6 generic map(INIT => "1111111011101100111011001100100011101100110010001100100010000000") port map( O =>C_1_S_4_out, I0 =>  C_1_S_4_L_0_out, I1 =>  C_1_S_4_L_1_out, I2 =>  C_1_S_4_L_2_out, I3 =>  C_1_S_4_L_3_out, I4 =>  C_1_S_4_L_4_out, I5 =>  C_1_S_4_L_5_out); 
C_1_S_5_inst : LUT6 generic map(INIT => "1111111111111110111111101100100011101100100000001000000000000000") port map( O =>C_1_S_5_out, I0 =>  C_1_S_5_L_0_out, I1 =>  C_1_S_5_L_1_out, I2 =>  C_1_S_5_L_2_out, I3 =>  C_1_S_5_L_3_out, I4 =>  C_1_S_5_L_4_out, I5 =>  C_1_S_5_L_5_out); 

C_1_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_1_out, I0 =>  C_1_S_0_out, I1 =>  C_1_S_1_out, I2 =>  C_1_S_2_out, I3 =>  C_1_S_3_out, I4 =>  C_1_S_4_out, I5 =>  C_1_S_5_out); 

 
C_2_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_2_S_0_out, I0 =>  C_2_S_0_L_0_out, I1 =>  C_2_S_0_L_1_out, I2 =>  C_2_S_0_L_2_out, I3 =>  C_2_S_0_L_3_out, I4 =>  C_2_S_0_L_4_out, I5 =>  C_2_S_0_L_5_out); 
C_2_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_2_S_1_out, I0 =>  C_2_S_1_L_0_out, I1 =>  C_2_S_1_L_1_out, I2 =>  C_2_S_1_L_2_out, I3 =>  C_2_S_1_L_3_out, I4 =>  C_2_S_1_L_4_out, I5 =>  C_2_S_1_L_5_out); 
C_2_S_2_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_2_S_2_out, I0 =>  C_2_S_2_L_0_out, I1 =>  C_2_S_2_L_1_out, I2 =>  C_2_S_2_L_2_out, I3 =>  C_2_S_2_L_3_out, I4 =>  C_2_S_2_L_4_out, I5 =>  C_2_S_2_L_5_out); 
C_2_S_3_inst : LUT6 generic map(INIT => "1111111011101000111111101110100011101000100000001110100010000000") port map( O =>C_2_S_3_out, I0 =>  C_2_S_3_L_0_out, I1 =>  C_2_S_3_L_1_out, I2 =>  C_2_S_3_L_2_out, I3 =>  C_2_S_3_L_3_out, I4 =>  C_2_S_3_L_4_out, I5 =>  C_2_S_3_L_5_out); 
C_2_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010001010100011101010111010001010100010000000") port map( O =>C_2_S_4_out, I0 =>  C_2_S_4_L_0_out, I1 =>  C_2_S_4_L_1_out, I2 =>  C_2_S_4_L_2_out, I3 =>  C_2_S_4_L_3_out, I4 =>  C_2_S_4_L_4_out, I5 =>  C_2_S_4_L_5_out); 
C_2_S_5_inst : LUT6 generic map(INIT => "1111111011101000111111101110100011101000100000001110100010000000") port map( O =>C_2_S_5_out, I0 =>  C_2_S_5_L_0_out, I1 =>  C_2_S_5_L_1_out, I2 =>  C_2_S_5_L_2_out, I3 =>  C_2_S_5_L_3_out, I4 =>  C_2_S_5_L_4_out, I5 =>  C_2_S_5_L_5_out); 

C_2_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_2_out, I0 =>  C_2_S_0_out, I1 =>  C_2_S_1_out, I2 =>  C_2_S_2_out, I3 =>  C_2_S_3_out, I4 =>  C_2_S_4_out, I5 =>  C_2_S_5_out); 

 
C_3_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_3_S_0_out, I0 =>  C_3_S_0_L_0_out, I1 =>  C_3_S_0_L_1_out, I2 =>  C_3_S_0_L_2_out, I3 =>  C_3_S_0_L_3_out, I4 =>  C_3_S_0_L_4_out, I5 =>  C_3_S_0_L_5_out); 
C_3_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_3_S_1_out, I0 =>  C_3_S_1_L_0_out, I1 =>  C_3_S_1_L_1_out, I2 =>  C_3_S_1_L_2_out, I3 =>  C_3_S_1_L_3_out, I4 =>  C_3_S_1_L_4_out, I5 =>  C_3_S_1_L_5_out); 
C_3_S_2_inst : LUT6 generic map(INIT => "1111111011111010111010001110100011101000111010001010000010000000") port map( O =>C_3_S_2_out, I0 =>  C_3_S_2_L_0_out, I1 =>  C_3_S_2_L_1_out, I2 =>  C_3_S_2_L_2_out, I3 =>  C_3_S_2_L_3_out, I4 =>  C_3_S_2_L_4_out, I5 =>  C_3_S_2_L_5_out); 
C_3_S_3_inst : LUT6 generic map(INIT => "1111111011111100111010001110100011101000111010001100000010000000") port map( O =>C_3_S_3_out, I0 =>  C_3_S_3_L_0_out, I1 =>  C_3_S_3_L_1_out, I2 =>  C_3_S_3_L_2_out, I3 =>  C_3_S_3_L_3_out, I4 =>  C_3_S_3_L_4_out, I5 =>  C_3_S_3_L_5_out); 
C_3_S_4_inst : LUT6 generic map(INIT => "1111111011101000111011001100100011101100110010001110100010000000") port map( O =>C_3_S_4_out, I0 =>  C_3_S_4_L_0_out, I1 =>  C_3_S_4_L_1_out, I2 =>  C_3_S_4_L_2_out, I3 =>  C_3_S_4_L_3_out, I4 =>  C_3_S_4_L_4_out, I5 =>  C_3_S_4_L_5_out); 
C_3_S_5_inst : LUT6 generic map(INIT => "1111111011111100111111001100000011111100110000001100000010000000") port map( O =>C_3_S_5_out, I0 =>  C_3_S_5_L_0_out, I1 =>  C_3_S_5_L_1_out, I2 =>  C_3_S_5_L_2_out, I3 =>  C_3_S_5_L_3_out, I4 =>  C_3_S_5_L_4_out, I5 =>  C_3_S_5_L_5_out); 

C_3_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_3_out, I0 =>  C_3_S_0_out, I1 =>  C_3_S_1_out, I2 =>  C_3_S_2_out, I3 =>  C_3_S_3_out, I4 =>  C_3_S_4_out, I5 =>  C_3_S_5_out); 

 
C_4_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_4_S_0_out, I0 =>  C_4_S_0_L_0_out, I1 =>  C_4_S_0_L_1_out, I2 =>  C_4_S_0_L_2_out, I3 =>  C_4_S_0_L_3_out, I4 =>  C_4_S_0_L_4_out, I5 =>  C_4_S_0_L_5_out); 
C_4_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_4_S_1_out, I0 =>  C_4_S_1_L_0_out, I1 =>  C_4_S_1_L_1_out, I2 =>  C_4_S_1_L_2_out, I3 =>  C_4_S_1_L_3_out, I4 =>  C_4_S_1_L_4_out, I5 =>  C_4_S_1_L_5_out); 
C_4_S_2_inst : LUT6 generic map(INIT => "1111111011101100111011001100100011101100110010001100100010000000") port map( O =>C_4_S_2_out, I0 =>  C_4_S_2_L_0_out, I1 =>  C_4_S_2_L_1_out, I2 =>  C_4_S_2_L_2_out, I3 =>  C_4_S_2_L_3_out, I4 =>  C_4_S_2_L_4_out, I5 =>  C_4_S_2_L_5_out); 
C_4_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001110100011101000111010001110100010000000") port map( O =>C_4_S_3_out, I0 =>  C_4_S_3_L_0_out, I1 =>  C_4_S_3_L_1_out, I2 =>  C_4_S_3_L_2_out, I3 =>  C_4_S_3_L_3_out, I4 =>  C_4_S_3_L_4_out, I5 =>  C_4_S_3_L_5_out); 
C_4_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_4_S_4_out, I0 =>  C_4_S_4_L_0_out, I1 =>  C_4_S_4_L_1_out, I2 =>  C_4_S_4_L_2_out, I3 =>  C_4_S_4_L_3_out, I4 =>  C_4_S_4_L_4_out, I5 =>  C_4_S_4_L_5_out); 
C_4_S_5_inst : LUT6 generic map(INIT => "1111111111111110111111101110100011101000100000001000000000000000") port map( O =>C_4_S_5_out, I0 =>  C_4_S_5_L_0_out, I1 =>  C_4_S_5_L_1_out, I2 =>  C_4_S_5_L_2_out, I3 =>  C_4_S_5_L_3_out, I4 =>  C_4_S_5_L_4_out, I5 =>  C_4_S_5_L_5_out); 

C_4_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_4_out, I0 =>  C_4_S_0_out, I1 =>  C_4_S_1_out, I2 =>  C_4_S_2_out, I3 =>  C_4_S_3_out, I4 =>  C_4_S_4_out, I5 =>  C_4_S_5_out); 

 
C_5_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_5_S_0_out, I0 =>  C_5_S_0_L_0_out, I1 =>  C_5_S_0_L_1_out, I2 =>  C_5_S_0_L_2_out, I3 =>  C_5_S_0_L_3_out, I4 =>  C_5_S_0_L_4_out, I5 =>  C_5_S_0_L_5_out); 
C_5_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101110100011101000101010001010100010000000") port map( O =>C_5_S_1_out, I0 =>  C_5_S_1_L_0_out, I1 =>  C_5_S_1_L_1_out, I2 =>  C_5_S_1_L_2_out, I3 =>  C_5_S_1_L_3_out, I4 =>  C_5_S_1_L_4_out, I5 =>  C_5_S_1_L_5_out); 
C_5_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001000100011101110111010001110100010000000") port map( O =>C_5_S_2_out, I0 =>  C_5_S_2_L_0_out, I1 =>  C_5_S_2_L_1_out, I2 =>  C_5_S_2_L_2_out, I3 =>  C_5_S_2_L_3_out, I4 =>  C_5_S_2_L_4_out, I5 =>  C_5_S_2_L_5_out); 
C_5_S_3_inst : LUT6 generic map(INIT => "1111111011111110111111001110100011101000110000001000000010000000") port map( O =>C_5_S_3_out, I0 =>  C_5_S_3_L_0_out, I1 =>  C_5_S_3_L_1_out, I2 =>  C_5_S_3_L_2_out, I3 =>  C_5_S_3_L_3_out, I4 =>  C_5_S_3_L_4_out, I5 =>  C_5_S_3_L_5_out); 
C_5_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010001000000011111110111010001010100010000000") port map( O =>C_5_S_4_out, I0 =>  C_5_S_4_L_0_out, I1 =>  C_5_S_4_L_1_out, I2 =>  C_5_S_4_L_2_out, I3 =>  C_5_S_4_L_3_out, I4 =>  C_5_S_4_L_4_out, I5 =>  C_5_S_4_L_5_out); 
C_5_S_5_inst : LUT6 generic map(INIT => "1111111111111110111111101110100011101000100000001000000000000000") port map( O =>C_5_S_5_out, I0 =>  C_5_S_5_L_0_out, I1 =>  C_5_S_5_L_1_out, I2 =>  C_5_S_5_L_2_out, I3 =>  C_5_S_5_L_3_out, I4 =>  C_5_S_5_L_4_out, I5 =>  C_5_S_5_L_5_out); 

C_5_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_5_out, I0 =>  C_5_S_0_out, I1 =>  C_5_S_1_out, I2 =>  C_5_S_2_out, I3 =>  C_5_S_3_out, I4 =>  C_5_S_4_out, I5 =>  C_5_S_5_out); 

 
C_6_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_6_S_0_out, I0 =>  C_6_S_0_L_0_out, I1 =>  C_6_S_0_L_1_out, I2 =>  C_6_S_0_L_2_out, I3 =>  C_6_S_0_L_3_out, I4 =>  C_6_S_0_L_4_out, I5 =>  C_6_S_0_L_5_out); 
C_6_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_6_S_1_out, I0 =>  C_6_S_1_L_0_out, I1 =>  C_6_S_1_L_1_out, I2 =>  C_6_S_1_L_2_out, I3 =>  C_6_S_1_L_3_out, I4 =>  C_6_S_1_L_4_out, I5 =>  C_6_S_1_L_5_out); 
C_6_S_2_inst : LUT6 generic map(INIT => "1111111011111010111110001110000011111000111000001010000010000000") port map( O =>C_6_S_2_out, I0 =>  C_6_S_2_L_0_out, I1 =>  C_6_S_2_L_1_out, I2 =>  C_6_S_2_L_2_out, I3 =>  C_6_S_2_L_3_out, I4 =>  C_6_S_2_L_4_out, I5 =>  C_6_S_2_L_5_out); 
C_6_S_3_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_6_S_3_out, I0 =>  C_6_S_3_L_0_out, I1 =>  C_6_S_3_L_1_out, I2 =>  C_6_S_3_L_2_out, I3 =>  C_6_S_3_L_3_out, I4 =>  C_6_S_3_L_4_out, I5 =>  C_6_S_3_L_5_out); 
C_6_S_4_inst : LUT6 generic map(INIT => "1111111011111110111010001110100011101000111010001000000010000000") port map( O =>C_6_S_4_out, I0 =>  C_6_S_4_L_0_out, I1 =>  C_6_S_4_L_1_out, I2 =>  C_6_S_4_L_2_out, I3 =>  C_6_S_4_L_3_out, I4 =>  C_6_S_4_L_4_out, I5 =>  C_6_S_4_L_5_out); 
C_6_S_5_inst : LUT6 generic map(INIT => "1111111011101000111110101010100011101010101000001110100010000000") port map( O =>C_6_S_5_out, I0 =>  C_6_S_5_L_0_out, I1 =>  C_6_S_5_L_1_out, I2 =>  C_6_S_5_L_2_out, I3 =>  C_6_S_5_L_3_out, I4 =>  C_6_S_5_L_4_out, I5 =>  C_6_S_5_L_5_out); 

C_6_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_6_out, I0 =>  C_6_S_0_out, I1 =>  C_6_S_1_out, I2 =>  C_6_S_2_out, I3 =>  C_6_S_3_out, I4 =>  C_6_S_4_out, I5 =>  C_6_S_5_out); 

 
C_7_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_7_S_0_out, I0 =>  C_7_S_0_L_0_out, I1 =>  C_7_S_0_L_1_out, I2 =>  C_7_S_0_L_2_out, I3 =>  C_7_S_0_L_3_out, I4 =>  C_7_S_0_L_4_out, I5 =>  C_7_S_0_L_5_out); 
C_7_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_7_S_1_out, I0 =>  C_7_S_1_L_0_out, I1 =>  C_7_S_1_L_1_out, I2 =>  C_7_S_1_L_2_out, I3 =>  C_7_S_1_L_3_out, I4 =>  C_7_S_1_L_4_out, I5 =>  C_7_S_1_L_5_out); 
C_7_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010001000000011111110111010001010100010000000") port map( O =>C_7_S_2_out, I0 =>  C_7_S_2_L_0_out, I1 =>  C_7_S_2_L_1_out, I2 =>  C_7_S_2_L_2_out, I3 =>  C_7_S_2_L_3_out, I4 =>  C_7_S_2_L_4_out, I5 =>  C_7_S_2_L_5_out); 
C_7_S_3_inst : LUT6 generic map(INIT => "1111111111111110111010001110100011101000111010001000000000000000") port map( O =>C_7_S_3_out, I0 =>  C_7_S_3_L_0_out, I1 =>  C_7_S_3_L_1_out, I2 =>  C_7_S_3_L_2_out, I3 =>  C_7_S_3_L_3_out, I4 =>  C_7_S_3_L_4_out, I5 =>  C_7_S_3_L_5_out); 
C_7_S_4_inst : LUT6 generic map(INIT => "1111111111101010111111101000000011111110100000001010100000000000") port map( O =>C_7_S_4_out, I0 =>  C_7_S_4_L_0_out, I1 =>  C_7_S_4_L_1_out, I2 =>  C_7_S_4_L_2_out, I3 =>  C_7_S_4_L_3_out, I4 =>  C_7_S_4_L_4_out, I5 =>  C_7_S_4_L_5_out); 
C_7_S_5_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_7_S_5_out, I0 =>  C_7_S_5_L_0_out, I1 =>  C_7_S_5_L_1_out, I2 =>  C_7_S_5_L_2_out, I3 =>  C_7_S_5_L_3_out, I4 =>  C_7_S_5_L_4_out, I5 =>  C_7_S_5_L_5_out); 

C_7_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_7_out, I0 =>  C_7_S_0_out, I1 =>  C_7_S_1_out, I2 =>  C_7_S_2_out, I3 =>  C_7_S_3_out, I4 =>  C_7_S_4_out, I5 =>  C_7_S_5_out); 

 
C_8_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_8_S_0_out, I0 =>  C_8_S_0_L_0_out, I1 =>  C_8_S_0_L_1_out, I2 =>  C_8_S_0_L_2_out, I3 =>  C_8_S_0_L_3_out, I4 =>  C_8_S_0_L_4_out, I5 =>  C_8_S_0_L_5_out); 
C_8_S_1_inst : LUT6 generic map(INIT => "1111101011101010101010101010100011101010101010101010100010100000") port map( O =>C_8_S_1_out, I0 =>  C_8_S_1_L_0_out, I1 =>  C_8_S_1_L_1_out, I2 =>  C_8_S_1_L_2_out, I3 =>  C_8_S_1_L_3_out, I4 =>  C_8_S_1_L_4_out, I5 =>  C_8_S_1_L_5_out); 
C_8_S_2_inst : LUT6 generic map(INIT => "1111111111101100111011001000000011111110110010001100100000000000") port map( O =>C_8_S_2_out, I0 =>  C_8_S_2_L_0_out, I1 =>  C_8_S_2_L_1_out, I2 =>  C_8_S_2_L_2_out, I3 =>  C_8_S_2_L_3_out, I4 =>  C_8_S_2_L_4_out, I5 =>  C_8_S_2_L_5_out); 
C_8_S_3_inst : LUT6 generic map(INIT => "1111111111111111111111101110100011101000100000000000000000000000") port map( O =>C_8_S_3_out, I0 =>  C_8_S_3_L_0_out, I1 =>  C_8_S_3_L_1_out, I2 =>  C_8_S_3_L_2_out, I3 =>  C_8_S_3_L_3_out, I4 =>  C_8_S_3_L_4_out, I5 =>  C_8_S_3_L_5_out); 
C_8_S_4_inst : LUT6 generic map(INIT => "1111111111101110111111101000000011111110100000001000100000000000") port map( O =>C_8_S_4_out, I0 =>  C_8_S_4_L_0_out, I1 =>  C_8_S_4_L_1_out, I2 =>  C_8_S_4_L_2_out, I3 =>  C_8_S_4_L_3_out, I4 =>  C_8_S_4_L_4_out, I5 =>  C_8_S_4_L_5_out); 
C_8_S_5_inst : LUT6 generic map(INIT => "1111111011111000111110101110100011101000101000001110000010000000") port map( O =>C_8_S_5_out, I0 =>  C_8_S_5_L_0_out, I1 =>  C_8_S_5_L_1_out, I2 =>  C_8_S_5_L_2_out, I3 =>  C_8_S_5_L_3_out, I4 =>  C_8_S_5_L_4_out, I5 =>  C_8_S_5_L_5_out); 

C_8_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_8_out, I0 =>  C_8_S_0_out, I1 =>  C_8_S_1_out, I2 =>  C_8_S_2_out, I3 =>  C_8_S_3_out, I4 =>  C_8_S_4_out, I5 =>  C_8_S_5_out); 

 
C_9_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_9_S_0_out, I0 =>  C_9_S_0_L_0_out, I1 =>  C_9_S_0_L_1_out, I2 =>  C_9_S_0_L_2_out, I3 =>  C_9_S_0_L_3_out, I4 =>  C_9_S_0_L_4_out, I5 =>  C_9_S_0_L_5_out); 
C_9_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_9_S_1_out, I0 =>  C_9_S_1_L_0_out, I1 =>  C_9_S_1_L_1_out, I2 =>  C_9_S_1_L_2_out, I3 =>  C_9_S_1_L_3_out, I4 =>  C_9_S_1_L_4_out, I5 =>  C_9_S_1_L_5_out); 
C_9_S_2_inst : LUT6 generic map(INIT => "1111111011101110111010001000100011101110111010001000100010000000") port map( O =>C_9_S_2_out, I0 =>  C_9_S_2_L_0_out, I1 =>  C_9_S_2_L_1_out, I2 =>  C_9_S_2_L_2_out, I3 =>  C_9_S_2_L_3_out, I4 =>  C_9_S_2_L_4_out, I5 =>  C_9_S_2_L_5_out); 
C_9_S_3_inst : LUT6 generic map(INIT => "1111111111111000111111101110000011111000100000001110000000000000") port map( O =>C_9_S_3_out, I0 =>  C_9_S_3_L_0_out, I1 =>  C_9_S_3_L_1_out, I2 =>  C_9_S_3_L_2_out, I3 =>  C_9_S_3_L_3_out, I4 =>  C_9_S_3_L_4_out, I5 =>  C_9_S_3_L_5_out); 
C_9_S_4_inst : LUT6 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_9_S_4_out, I0 =>  C_9_S_4_L_0_out, I1 =>  C_9_S_4_L_1_out, I2 =>  C_9_S_4_L_2_out, I3 =>  C_9_S_4_L_3_out, I4 =>  C_9_S_4_L_4_out, I5 =>  C_9_S_4_L_5_out); 
C_9_S_5_inst : LUT6 generic map(INIT => "1111111111101100111011001000000011111110110010001100100000000000") port map( O =>C_9_S_5_out, I0 =>  C_9_S_5_L_0_out, I1 =>  C_9_S_5_L_1_out, I2 =>  C_9_S_5_L_2_out, I3 =>  C_9_S_5_L_3_out, I4 =>  C_9_S_5_L_4_out, I5 =>  C_9_S_5_L_5_out); 

C_9_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_9_out, I0 =>  C_9_S_0_out, I1 =>  C_9_S_1_out, I2 =>  C_9_S_2_out, I3 =>  C_9_S_3_out, I4 =>  C_9_S_4_out, I5 =>  C_9_S_5_out); 

 
C_10_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_10_S_0_out, I0 =>  C_10_S_0_L_0_out, I1 =>  C_10_S_0_L_1_out, I2 =>  C_10_S_0_L_2_out, I3 =>  C_10_S_0_L_3_out, I4 =>  C_10_S_0_L_4_out, I5 =>  C_10_S_0_L_5_out); 
C_10_S_1_inst : LUT6 generic map(INIT => "1111111011101000111011101110100011101000100010001110100010000000") port map( O =>C_10_S_1_out, I0 =>  C_10_S_1_L_0_out, I1 =>  C_10_S_1_L_1_out, I2 =>  C_10_S_1_L_2_out, I3 =>  C_10_S_1_L_3_out, I4 =>  C_10_S_1_L_4_out, I5 =>  C_10_S_1_L_5_out); 
C_10_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_10_S_2_out, I0 =>  C_10_S_2_L_0_out, I1 =>  C_10_S_2_L_1_out, I2 =>  C_10_S_2_L_2_out, I3 =>  C_10_S_2_L_3_out, I4 =>  C_10_S_2_L_4_out, I5 =>  C_10_S_2_L_5_out); 
C_10_S_3_inst : LUT6 generic map(INIT => "1111111011101100111011001100100011101100110010001100100010000000") port map( O =>C_10_S_3_out, I0 =>  C_10_S_3_L_0_out, I1 =>  C_10_S_3_L_1_out, I2 =>  C_10_S_3_L_2_out, I3 =>  C_10_S_3_L_3_out, I4 =>  C_10_S_3_L_4_out, I5 =>  C_10_S_3_L_5_out); 
C_10_S_4_inst : LUT6 generic map(INIT => "1111111011101000111011101000100011101110100010001110100010000000") port map( O =>C_10_S_4_out, I0 =>  C_10_S_4_L_0_out, I1 =>  C_10_S_4_L_1_out, I2 =>  C_10_S_4_L_2_out, I3 =>  C_10_S_4_L_3_out, I4 =>  C_10_S_4_L_4_out, I5 =>  C_10_S_4_L_5_out); 
C_10_S_5_inst : LUT6 generic map(INIT => "1111111111101010111111101010100011101010100000001010100000000000") port map( O =>C_10_S_5_out, I0 =>  C_10_S_5_L_0_out, I1 =>  C_10_S_5_L_1_out, I2 =>  C_10_S_5_L_2_out, I3 =>  C_10_S_5_L_3_out, I4 =>  C_10_S_5_L_4_out, I5 =>  C_10_S_5_L_5_out); 

C_10_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_10_out, I0 =>  C_10_S_0_out, I1 =>  C_10_S_1_out, I2 =>  C_10_S_2_out, I3 =>  C_10_S_3_out, I4 =>  C_10_S_4_out, I5 =>  C_10_S_5_out); 

 
C_11_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_11_S_0_out, I0 =>  C_11_S_0_L_0_out, I1 =>  C_11_S_0_L_1_out, I2 =>  C_11_S_0_L_2_out, I3 =>  C_11_S_0_L_3_out, I4 =>  C_11_S_0_L_4_out, I5 =>  C_11_S_0_L_5_out); 
C_11_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010101010100011101010101010001110100010000000") port map( O =>C_11_S_1_out, I0 =>  C_11_S_1_L_0_out, I1 =>  C_11_S_1_L_1_out, I2 =>  C_11_S_1_L_2_out, I3 =>  C_11_S_1_L_3_out, I4 =>  C_11_S_1_L_4_out, I5 =>  C_11_S_1_L_5_out); 
C_11_S_2_inst : LUT6 generic map(INIT => "1111111111101000111010101000000011111110101010001110100000000000") port map( O =>C_11_S_2_out, I0 =>  C_11_S_2_L_0_out, I1 =>  C_11_S_2_L_1_out, I2 =>  C_11_S_2_L_2_out, I3 =>  C_11_S_2_L_3_out, I4 =>  C_11_S_2_L_4_out, I5 =>  C_11_S_2_L_5_out); 
C_11_S_3_inst : LUT6 generic map(INIT => "1111111111111110111111101110100011101000100000001000000000000000") port map( O =>C_11_S_3_out, I0 =>  C_11_S_3_L_0_out, I1 =>  C_11_S_3_L_1_out, I2 =>  C_11_S_3_L_2_out, I3 =>  C_11_S_3_L_3_out, I4 =>  C_11_S_3_L_4_out, I5 =>  C_11_S_3_L_5_out); 
C_11_S_4_inst : LUT6 generic map(INIT => "1111111011101010111111101010100011101010100000001010100010000000") port map( O =>C_11_S_4_out, I0 =>  C_11_S_4_L_0_out, I1 =>  C_11_S_4_L_1_out, I2 =>  C_11_S_4_L_2_out, I3 =>  C_11_S_4_L_3_out, I4 =>  C_11_S_4_L_4_out, I5 =>  C_11_S_4_L_5_out); 
C_11_S_5_inst : LUT6 generic map(INIT => "1111111111101100111011001000000011111110110010001100100000000000") port map( O =>C_11_S_5_out, I0 =>  C_11_S_5_L_0_out, I1 =>  C_11_S_5_L_1_out, I2 =>  C_11_S_5_L_2_out, I3 =>  C_11_S_5_L_3_out, I4 =>  C_11_S_5_L_4_out, I5 =>  C_11_S_5_L_5_out); 

C_11_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_11_out, I0 =>  C_11_S_0_out, I1 =>  C_11_S_1_out, I2 =>  C_11_S_2_out, I3 =>  C_11_S_3_out, I4 =>  C_11_S_4_out, I5 =>  C_11_S_5_out); 

 
C_12_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_12_S_0_out, I0 =>  C_12_S_0_L_0_out, I1 =>  C_12_S_0_L_1_out, I2 =>  C_12_S_0_L_2_out, I3 =>  C_12_S_0_L_3_out, I4 =>  C_12_S_0_L_4_out, I5 =>  C_12_S_0_L_5_out); 
C_12_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_12_S_1_out, I0 =>  C_12_S_1_L_0_out, I1 =>  C_12_S_1_L_1_out, I2 =>  C_12_S_1_L_2_out, I3 =>  C_12_S_1_L_3_out, I4 =>  C_12_S_1_L_4_out, I5 =>  C_12_S_1_L_5_out); 
C_12_S_2_inst : LUT6 generic map(INIT => "1111111011101100111011001100100011101100110010001100100010000000") port map( O =>C_12_S_2_out, I0 =>  C_12_S_2_L_0_out, I1 =>  C_12_S_2_L_1_out, I2 =>  C_12_S_2_L_2_out, I3 =>  C_12_S_2_L_3_out, I4 =>  C_12_S_2_L_4_out, I5 =>  C_12_S_2_L_5_out); 
C_12_S_3_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_12_S_3_out, I0 =>  C_12_S_3_L_0_out, I1 =>  C_12_S_3_L_1_out, I2 =>  C_12_S_3_L_2_out, I3 =>  C_12_S_3_L_3_out, I4 =>  C_12_S_3_L_4_out, I5 =>  C_12_S_3_L_5_out); 
C_12_S_4_inst : LUT6 generic map(INIT => "1111111111101100111011101100100011101100100010001100100000000000") port map( O =>C_12_S_4_out, I0 =>  C_12_S_4_L_0_out, I1 =>  C_12_S_4_L_1_out, I2 =>  C_12_S_4_L_2_out, I3 =>  C_12_S_4_L_3_out, I4 =>  C_12_S_4_L_4_out, I5 =>  C_12_S_4_L_5_out); 
C_12_S_5_inst : LUT6 generic map(INIT => "1111111111111100111111001100000011111100110000001100000000000000") port map( O =>C_12_S_5_out, I0 =>  C_12_S_5_L_0_out, I1 =>  C_12_S_5_L_1_out, I2 =>  C_12_S_5_L_2_out, I3 =>  C_12_S_5_L_3_out, I4 =>  C_12_S_5_L_4_out, I5 =>  C_12_S_5_L_5_out); 

C_12_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_12_out, I0 =>  C_12_S_0_out, I1 =>  C_12_S_1_out, I2 =>  C_12_S_2_out, I3 =>  C_12_S_3_out, I4 =>  C_12_S_4_out, I5 =>  C_12_S_5_out); 

 
C_13_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_13_S_0_out, I0 =>  C_13_S_0_L_0_out, I1 =>  C_13_S_0_L_1_out, I2 =>  C_13_S_0_L_2_out, I3 =>  C_13_S_0_L_3_out, I4 =>  C_13_S_0_L_4_out, I5 =>  C_13_S_0_L_5_out); 
C_13_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010001110100011101000111010001110100010000000") port map( O =>C_13_S_1_out, I0 =>  C_13_S_1_L_0_out, I1 =>  C_13_S_1_L_1_out, I2 =>  C_13_S_1_L_2_out, I3 =>  C_13_S_1_L_3_out, I4 =>  C_13_S_1_L_4_out, I5 =>  C_13_S_1_L_5_out); 
C_13_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_13_S_2_out, I0 =>  C_13_S_2_L_0_out, I1 =>  C_13_S_2_L_1_out, I2 =>  C_13_S_2_L_2_out, I3 =>  C_13_S_2_L_3_out, I4 =>  C_13_S_2_L_4_out, I5 =>  C_13_S_2_L_5_out); 
C_13_S_3_inst : LUT6 generic map(INIT => "1111111111101010111010101000100011101110101010001010100000000000") port map( O =>C_13_S_3_out, I0 =>  C_13_S_3_L_0_out, I1 =>  C_13_S_3_L_1_out, I2 =>  C_13_S_3_L_2_out, I3 =>  C_13_S_3_L_3_out, I4 =>  C_13_S_3_L_4_out, I5 =>  C_13_S_3_L_5_out); 
C_13_S_4_inst : LUT6 generic map(INIT => "1111111111111100111111001110100011101000110000001100000000000000") port map( O =>C_13_S_4_out, I0 =>  C_13_S_4_L_0_out, I1 =>  C_13_S_4_L_1_out, I2 =>  C_13_S_4_L_2_out, I3 =>  C_13_S_4_L_3_out, I4 =>  C_13_S_4_L_4_out, I5 =>  C_13_S_4_L_5_out); 
C_13_S_5_inst : LUT6 generic map(INIT => "1111111011101100111011001100100011101100110010001100100010000000") port map( O =>C_13_S_5_out, I0 =>  C_13_S_5_L_0_out, I1 =>  C_13_S_5_L_1_out, I2 =>  C_13_S_5_L_2_out, I3 =>  C_13_S_5_L_3_out, I4 =>  C_13_S_5_L_4_out, I5 =>  C_13_S_5_L_5_out); 

C_13_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_13_out, I0 =>  C_13_S_0_out, I1 =>  C_13_S_1_out, I2 =>  C_13_S_2_out, I3 =>  C_13_S_3_out, I4 =>  C_13_S_4_out, I5 =>  C_13_S_5_out); 

 
C_14_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_14_S_0_out, I0 =>  C_14_S_0_L_0_out, I1 =>  C_14_S_0_L_1_out, I2 =>  C_14_S_0_L_2_out, I3 =>  C_14_S_0_L_3_out, I4 =>  C_14_S_0_L_4_out, I5 =>  C_14_S_0_L_5_out); 
C_14_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101110100011101000101010001010100010000000") port map( O =>C_14_S_1_out, I0 =>  C_14_S_1_L_0_out, I1 =>  C_14_S_1_L_1_out, I2 =>  C_14_S_1_L_2_out, I3 =>  C_14_S_1_L_3_out, I4 =>  C_14_S_1_L_4_out, I5 =>  C_14_S_1_L_5_out); 
C_14_S_2_inst : LUT6 generic map(INIT => "1111111111101110111111101100100011101100100000001000100000000000") port map( O =>C_14_S_2_out, I0 =>  C_14_S_2_L_0_out, I1 =>  C_14_S_2_L_1_out, I2 =>  C_14_S_2_L_2_out, I3 =>  C_14_S_2_L_3_out, I4 =>  C_14_S_2_L_4_out, I5 =>  C_14_S_2_L_5_out); 
C_14_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001100100011101100111010001110100010000000") port map( O =>C_14_S_3_out, I0 =>  C_14_S_3_L_0_out, I1 =>  C_14_S_3_L_1_out, I2 =>  C_14_S_3_L_2_out, I3 =>  C_14_S_3_L_3_out, I4 =>  C_14_S_3_L_4_out, I5 =>  C_14_S_3_L_5_out); 
C_14_S_4_inst : LUT6 generic map(INIT => "1111111111101010111010101000000011111110101010001010100000000000") port map( O =>C_14_S_4_out, I0 =>  C_14_S_4_L_0_out, I1 =>  C_14_S_4_L_1_out, I2 =>  C_14_S_4_L_2_out, I3 =>  C_14_S_4_L_3_out, I4 =>  C_14_S_4_L_4_out, I5 =>  C_14_S_4_L_5_out); 
C_14_S_5_inst : LUT6 generic map(INIT => "1111111111111100111111001100000011111100110000001100000000000000") port map( O =>C_14_S_5_out, I0 =>  C_14_S_5_L_0_out, I1 =>  C_14_S_5_L_1_out, I2 =>  C_14_S_5_L_2_out, I3 =>  C_14_S_5_L_3_out, I4 =>  C_14_S_5_L_4_out, I5 =>  C_14_S_5_L_5_out); 

C_14_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_14_out, I0 =>  C_14_S_0_out, I1 =>  C_14_S_1_out, I2 =>  C_14_S_2_out, I3 =>  C_14_S_3_out, I4 =>  C_14_S_4_out, I5 =>  C_14_S_5_out); 

 
C_15_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_15_S_0_out, I0 =>  C_15_S_0_L_0_out, I1 =>  C_15_S_0_L_1_out, I2 =>  C_15_S_0_L_2_out, I3 =>  C_15_S_0_L_3_out, I4 =>  C_15_S_0_L_4_out, I5 =>  C_15_S_0_L_5_out); 
C_15_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101110100011101000101010001010100010000000") port map( O =>C_15_S_1_out, I0 =>  C_15_S_1_L_0_out, I1 =>  C_15_S_1_L_1_out, I2 =>  C_15_S_1_L_2_out, I3 =>  C_15_S_1_L_3_out, I4 =>  C_15_S_1_L_4_out, I5 =>  C_15_S_1_L_5_out); 
C_15_S_2_inst : LUT6 generic map(INIT => "1111111111111110111010101010000011111010101010001000000000000000") port map( O =>C_15_S_2_out, I0 =>  C_15_S_2_L_0_out, I1 =>  C_15_S_2_L_1_out, I2 =>  C_15_S_2_L_2_out, I3 =>  C_15_S_2_L_3_out, I4 =>  C_15_S_2_L_4_out, I5 =>  C_15_S_2_L_5_out); 
C_15_S_3_inst : LUT6 generic map(INIT => "1111111011101010111010101000100011101110101010001010100010000000") port map( O =>C_15_S_3_out, I0 =>  C_15_S_3_L_0_out, I1 =>  C_15_S_3_L_1_out, I2 =>  C_15_S_3_L_2_out, I3 =>  C_15_S_3_L_3_out, I4 =>  C_15_S_3_L_4_out, I5 =>  C_15_S_3_L_5_out); 
C_15_S_4_inst : LUT6 generic map(INIT => "1111111111111000111110001000000011111110111000001110000000000000") port map( O =>C_15_S_4_out, I0 =>  C_15_S_4_L_0_out, I1 =>  C_15_S_4_L_1_out, I2 =>  C_15_S_4_L_2_out, I3 =>  C_15_S_4_L_3_out, I4 =>  C_15_S_4_L_4_out, I5 =>  C_15_S_4_L_5_out); 
C_15_S_5_inst : LUT6 generic map(INIT => "1111111111111000111111001110000011111000110000001110000000000000") port map( O =>C_15_S_5_out, I0 =>  C_15_S_5_L_0_out, I1 =>  C_15_S_5_L_1_out, I2 =>  C_15_S_5_L_2_out, I3 =>  C_15_S_5_L_3_out, I4 =>  C_15_S_5_L_4_out, I5 =>  C_15_S_5_L_5_out); 

C_15_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_15_out, I0 =>  C_15_S_0_out, I1 =>  C_15_S_1_out, I2 =>  C_15_S_2_out, I3 =>  C_15_S_3_out, I4 =>  C_15_S_4_out, I5 =>  C_15_S_5_out); 

 
C_16_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_16_S_0_out, I0 =>  C_16_S_0_L_0_out, I1 =>  C_16_S_0_L_1_out, I2 =>  C_16_S_0_L_2_out, I3 =>  C_16_S_0_L_3_out, I4 =>  C_16_S_0_L_4_out, I5 =>  C_16_S_0_L_5_out); 
C_16_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_16_S_1_out, I0 =>  C_16_S_1_L_0_out, I1 =>  C_16_S_1_L_1_out, I2 =>  C_16_S_1_L_2_out, I3 =>  C_16_S_1_L_3_out, I4 =>  C_16_S_1_L_4_out, I5 =>  C_16_S_1_L_5_out); 
C_16_S_2_inst : LUT6 generic map(INIT => "1111111111101100111011001100100011101100110010001100100000000000") port map( O =>C_16_S_2_out, I0 =>  C_16_S_2_L_0_out, I1 =>  C_16_S_2_L_1_out, I2 =>  C_16_S_2_L_2_out, I3 =>  C_16_S_2_L_3_out, I4 =>  C_16_S_2_L_4_out, I5 =>  C_16_S_2_L_5_out); 
C_16_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_16_S_3_out, I0 =>  C_16_S_3_L_0_out, I1 =>  C_16_S_3_L_1_out, I2 =>  C_16_S_3_L_2_out, I3 =>  C_16_S_3_L_3_out, I4 =>  C_16_S_3_L_4_out, I5 =>  C_16_S_3_L_5_out); 
C_16_S_4_inst : LUT6 generic map(INIT => "1111111111111100111111001100000011111100110000001100000000000000") port map( O =>C_16_S_4_out, I0 =>  C_16_S_4_L_0_out, I1 =>  C_16_S_4_L_1_out, I2 =>  C_16_S_4_L_2_out, I3 =>  C_16_S_4_L_3_out, I4 =>  C_16_S_4_L_4_out, I5 =>  C_16_S_4_L_5_out); 
C_16_S_5_inst : LUT6 generic map(INIT => "1111111011101010111010101010000011111010101010001010100010000000") port map( O =>C_16_S_5_out, I0 =>  C_16_S_5_L_0_out, I1 =>  C_16_S_5_L_1_out, I2 =>  C_16_S_5_L_2_out, I3 =>  C_16_S_5_L_3_out, I4 =>  C_16_S_5_L_4_out, I5 =>  C_16_S_5_L_5_out); 

C_16_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_16_out, I0 =>  C_16_S_0_out, I1 =>  C_16_S_1_out, I2 =>  C_16_S_2_out, I3 =>  C_16_S_3_out, I4 =>  C_16_S_4_out, I5 =>  C_16_S_5_out); 

 
C_17_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_17_S_0_out, I0 =>  C_17_S_0_L_0_out, I1 =>  C_17_S_0_L_1_out, I2 =>  C_17_S_0_L_2_out, I3 =>  C_17_S_0_L_3_out, I4 =>  C_17_S_0_L_4_out, I5 =>  C_17_S_0_L_5_out); 
C_17_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_17_S_1_out, I0 =>  C_17_S_1_L_0_out, I1 =>  C_17_S_1_L_1_out, I2 =>  C_17_S_1_L_2_out, I3 =>  C_17_S_1_L_3_out, I4 =>  C_17_S_1_L_4_out, I5 =>  C_17_S_1_L_5_out); 
C_17_S_2_inst : LUT6 generic map(INIT => "1111111011111100111111001110100011101000110000001100000010000000") port map( O =>C_17_S_2_out, I0 =>  C_17_S_2_L_0_out, I1 =>  C_17_S_2_L_1_out, I2 =>  C_17_S_2_L_2_out, I3 =>  C_17_S_2_L_3_out, I4 =>  C_17_S_2_L_4_out, I5 =>  C_17_S_2_L_5_out); 
C_17_S_3_inst : LUT6 generic map(INIT => "1111111111111110111110101110100011101000101000001000000000000000") port map( O =>C_17_S_3_out, I0 =>  C_17_S_3_L_0_out, I1 =>  C_17_S_3_L_1_out, I2 =>  C_17_S_3_L_2_out, I3 =>  C_17_S_3_L_3_out, I4 =>  C_17_S_3_L_4_out, I5 =>  C_17_S_3_L_5_out); 
C_17_S_4_inst : LUT6 generic map(INIT => "1111111111111010111110101010000011111010101000001010000000000000") port map( O =>C_17_S_4_out, I0 =>  C_17_S_4_L_0_out, I1 =>  C_17_S_4_L_1_out, I2 =>  C_17_S_4_L_2_out, I3 =>  C_17_S_4_L_3_out, I4 =>  C_17_S_4_L_4_out, I5 =>  C_17_S_4_L_5_out); 
C_17_S_5_inst : LUT6 generic map(INIT => "1111111111101000111011101000100011101110100010001110100000000000") port map( O =>C_17_S_5_out, I0 =>  C_17_S_5_L_0_out, I1 =>  C_17_S_5_L_1_out, I2 =>  C_17_S_5_L_2_out, I3 =>  C_17_S_5_L_3_out, I4 =>  C_17_S_5_L_4_out, I5 =>  C_17_S_5_L_5_out); 

C_17_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_17_out, I0 =>  C_17_S_0_out, I1 =>  C_17_S_1_out, I2 =>  C_17_S_2_out, I3 =>  C_17_S_3_out, I4 =>  C_17_S_4_out, I5 =>  C_17_S_5_out); 

 
C_18_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_18_S_0_out, I0 =>  C_18_S_0_L_0_out, I1 =>  C_18_S_0_L_1_out, I2 =>  C_18_S_0_L_2_out, I3 =>  C_18_S_0_L_3_out, I4 =>  C_18_S_0_L_4_out, I5 =>  C_18_S_0_L_5_out); 
C_18_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_18_S_1_out, I0 =>  C_18_S_1_L_0_out, I1 =>  C_18_S_1_L_1_out, I2 =>  C_18_S_1_L_2_out, I3 =>  C_18_S_1_L_3_out, I4 =>  C_18_S_1_L_4_out, I5 =>  C_18_S_1_L_5_out); 
C_18_S_2_inst : LUT6 generic map(INIT => "1111111111111110111010001000000011111110111010001000000000000000") port map( O =>C_18_S_2_out, I0 =>  C_18_S_2_L_0_out, I1 =>  C_18_S_2_L_1_out, I2 =>  C_18_S_2_L_2_out, I3 =>  C_18_S_2_L_3_out, I4 =>  C_18_S_2_L_4_out, I5 =>  C_18_S_2_L_5_out); 
C_18_S_3_inst : LUT6 generic map(INIT => "1111111011101110111010101010100011101010101010001000100010000000") port map( O =>C_18_S_3_out, I0 =>  C_18_S_3_L_0_out, I1 =>  C_18_S_3_L_1_out, I2 =>  C_18_S_3_L_2_out, I3 =>  C_18_S_3_L_3_out, I4 =>  C_18_S_3_L_4_out, I5 =>  C_18_S_3_L_5_out); 
C_18_S_4_inst : LUT6 generic map(INIT => "1111111011111010111010101010100011101010101010001010000010000000") port map( O =>C_18_S_4_out, I0 =>  C_18_S_4_L_0_out, I1 =>  C_18_S_4_L_1_out, I2 =>  C_18_S_4_L_2_out, I3 =>  C_18_S_4_L_3_out, I4 =>  C_18_S_4_L_4_out, I5 =>  C_18_S_4_L_5_out); 
C_18_S_5_inst : LUT6 generic map(INIT => "1111111111111110111010101000000011111110101010001000000000000000") port map( O =>C_18_S_5_out, I0 =>  C_18_S_5_L_0_out, I1 =>  C_18_S_5_L_1_out, I2 =>  C_18_S_5_L_2_out, I3 =>  C_18_S_5_L_3_out, I4 =>  C_18_S_5_L_4_out, I5 =>  C_18_S_5_L_5_out); 

C_18_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_18_out, I0 =>  C_18_S_0_out, I1 =>  C_18_S_1_out, I2 =>  C_18_S_2_out, I3 =>  C_18_S_3_out, I4 =>  C_18_S_4_out, I5 =>  C_18_S_5_out); 

 
C_19_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_19_S_0_out, I0 =>  C_19_S_0_L_0_out, I1 =>  C_19_S_0_L_1_out, I2 =>  C_19_S_0_L_2_out, I3 =>  C_19_S_0_L_3_out, I4 =>  C_19_S_0_L_4_out, I5 =>  C_19_S_0_L_5_out); 
C_19_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_19_S_1_out, I0 =>  C_19_S_1_L_0_out, I1 =>  C_19_S_1_L_1_out, I2 =>  C_19_S_1_L_2_out, I3 =>  C_19_S_1_L_3_out, I4 =>  C_19_S_1_L_4_out, I5 =>  C_19_S_1_L_5_out); 
C_19_S_2_inst : LUT6 generic map(INIT => "1111111011101000111111001100000011111100110000001110100010000000") port map( O =>C_19_S_2_out, I0 =>  C_19_S_2_L_0_out, I1 =>  C_19_S_2_L_1_out, I2 =>  C_19_S_2_L_2_out, I3 =>  C_19_S_2_L_3_out, I4 =>  C_19_S_2_L_4_out, I5 =>  C_19_S_2_L_5_out); 
C_19_S_3_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_19_S_3_out, I0 =>  C_19_S_3_L_0_out, I1 =>  C_19_S_3_L_1_out, I2 =>  C_19_S_3_L_2_out, I3 =>  C_19_S_3_L_3_out, I4 =>  C_19_S_3_L_4_out, I5 =>  C_19_S_3_L_5_out); 
C_19_S_4_inst : LUT6 generic map(INIT => "1111111111111000111110001100000011111100111000001110000000000000") port map( O =>C_19_S_4_out, I0 =>  C_19_S_4_L_0_out, I1 =>  C_19_S_4_L_1_out, I2 =>  C_19_S_4_L_2_out, I3 =>  C_19_S_4_L_3_out, I4 =>  C_19_S_4_L_4_out, I5 =>  C_19_S_4_L_5_out); 
C_19_S_5_inst : LUT6 generic map(INIT => "1111111111111110111111101110000011111000100000001000000000000000") port map( O =>C_19_S_5_out, I0 =>  C_19_S_5_L_0_out, I1 =>  C_19_S_5_L_1_out, I2 =>  C_19_S_5_L_2_out, I3 =>  C_19_S_5_L_3_out, I4 =>  C_19_S_5_L_4_out, I5 =>  C_19_S_5_L_5_out); 

C_19_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_19_out, I0 =>  C_19_S_0_out, I1 =>  C_19_S_1_out, I2 =>  C_19_S_2_out, I3 =>  C_19_S_3_out, I4 =>  C_19_S_4_out, I5 =>  C_19_S_5_out); 

 
C_20_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_20_S_0_out, I0 =>  C_20_S_0_L_0_out, I1 =>  C_20_S_0_L_1_out, I2 =>  C_20_S_0_L_2_out, I3 =>  C_20_S_0_L_3_out, I4 =>  C_20_S_0_L_4_out, I5 =>  C_20_S_0_L_5_out); 
C_20_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010101110100011101000101010001110100010000000") port map( O =>C_20_S_1_out, I0 =>  C_20_S_1_L_0_out, I1 =>  C_20_S_1_L_1_out, I2 =>  C_20_S_1_L_2_out, I3 =>  C_20_S_1_L_3_out, I4 =>  C_20_S_1_L_4_out, I5 =>  C_20_S_1_L_5_out); 
C_20_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010101010100011101010101010001110100010000000") port map( O =>C_20_S_2_out, I0 =>  C_20_S_2_L_0_out, I1 =>  C_20_S_2_L_1_out, I2 =>  C_20_S_2_L_2_out, I3 =>  C_20_S_2_L_3_out, I4 =>  C_20_S_2_L_4_out, I5 =>  C_20_S_2_L_5_out); 
C_20_S_3_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_20_S_3_out, I0 =>  C_20_S_3_L_0_out, I1 =>  C_20_S_3_L_1_out, I2 =>  C_20_S_3_L_2_out, I3 =>  C_20_S_3_L_3_out, I4 =>  C_20_S_3_L_4_out, I5 =>  C_20_S_3_L_5_out); 
C_20_S_4_inst : LUT6 generic map(INIT => "1111111011101000111010001100100011101100111010001110100010000000") port map( O =>C_20_S_4_out, I0 =>  C_20_S_4_L_0_out, I1 =>  C_20_S_4_L_1_out, I2 =>  C_20_S_4_L_2_out, I3 =>  C_20_S_4_L_3_out, I4 =>  C_20_S_4_L_4_out, I5 =>  C_20_S_4_L_5_out); 
C_20_S_5_inst : LUT6 generic map(INIT => "1111111111111110111111001000000011111110110000001000000000000000") port map( O =>C_20_S_5_out, I0 =>  C_20_S_5_L_0_out, I1 =>  C_20_S_5_L_1_out, I2 =>  C_20_S_5_L_2_out, I3 =>  C_20_S_5_L_3_out, I4 =>  C_20_S_5_L_4_out, I5 =>  C_20_S_5_L_5_out); 

C_20_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_20_out, I0 =>  C_20_S_0_out, I1 =>  C_20_S_1_out, I2 =>  C_20_S_2_out, I3 =>  C_20_S_3_out, I4 =>  C_20_S_4_out, I5 =>  C_20_S_5_out); 

 
C_21_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_21_S_0_out, I0 =>  C_21_S_0_L_0_out, I1 =>  C_21_S_0_L_1_out, I2 =>  C_21_S_0_L_2_out, I3 =>  C_21_S_0_L_3_out, I4 =>  C_21_S_0_L_4_out, I5 =>  C_21_S_0_L_5_out); 
C_21_S_1_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_21_S_1_out, I0 =>  C_21_S_1_L_0_out, I1 =>  C_21_S_1_L_1_out, I2 =>  C_21_S_1_L_2_out, I3 =>  C_21_S_1_L_3_out, I4 =>  C_21_S_1_L_4_out, I5 =>  C_21_S_1_L_5_out); 
C_21_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_21_S_2_out, I0 =>  C_21_S_2_L_0_out, I1 =>  C_21_S_2_L_1_out, I2 =>  C_21_S_2_L_2_out, I3 =>  C_21_S_2_L_3_out, I4 =>  C_21_S_2_L_4_out, I5 =>  C_21_S_2_L_5_out); 
C_21_S_3_inst : LUT6 generic map(INIT => "1111111111101100111010001000000011111110111010001100100000000000") port map( O =>C_21_S_3_out, I0 =>  C_21_S_3_L_0_out, I1 =>  C_21_S_3_L_1_out, I2 =>  C_21_S_3_L_2_out, I3 =>  C_21_S_3_L_3_out, I4 =>  C_21_S_3_L_4_out, I5 =>  C_21_S_3_L_5_out); 
C_21_S_4_inst : LUT6 generic map(INIT => "1111111111111110111111001110100011101000110000001000000000000000") port map( O =>C_21_S_4_out, I0 =>  C_21_S_4_L_0_out, I1 =>  C_21_S_4_L_1_out, I2 =>  C_21_S_4_L_2_out, I3 =>  C_21_S_4_L_3_out, I4 =>  C_21_S_4_L_4_out, I5 =>  C_21_S_4_L_5_out); 
C_21_S_5_inst : LUT6 generic map(INIT => "1111111011111110111010101010100011101010101010001000000010000000") port map( O =>C_21_S_5_out, I0 =>  C_21_S_5_L_0_out, I1 =>  C_21_S_5_L_1_out, I2 =>  C_21_S_5_L_2_out, I3 =>  C_21_S_5_L_3_out, I4 =>  C_21_S_5_L_4_out, I5 =>  C_21_S_5_L_5_out); 

C_21_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_21_out, I0 =>  C_21_S_0_out, I1 =>  C_21_S_1_out, I2 =>  C_21_S_2_out, I3 =>  C_21_S_3_out, I4 =>  C_21_S_4_out, I5 =>  C_21_S_5_out); 

 
C_22_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_22_S_0_out, I0 =>  C_22_S_0_L_0_out, I1 =>  C_22_S_0_L_1_out, I2 =>  C_22_S_0_L_2_out, I3 =>  C_22_S_0_L_3_out, I4 =>  C_22_S_0_L_4_out, I5 =>  C_22_S_0_L_5_out); 
C_22_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_22_S_1_out, I0 =>  C_22_S_1_L_0_out, I1 =>  C_22_S_1_L_1_out, I2 =>  C_22_S_1_L_2_out, I3 =>  C_22_S_1_L_3_out, I4 =>  C_22_S_1_L_4_out, I5 =>  C_22_S_1_L_5_out); 
C_22_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001000100011101110111010001110100010000000") port map( O =>C_22_S_2_out, I0 =>  C_22_S_2_L_0_out, I1 =>  C_22_S_2_L_1_out, I2 =>  C_22_S_2_L_2_out, I3 =>  C_22_S_2_L_3_out, I4 =>  C_22_S_2_L_4_out, I5 =>  C_22_S_2_L_5_out); 
C_22_S_3_inst : LUT6 generic map(INIT => "1111111011111110111111101110100011101000100000001000000010000000") port map( O =>C_22_S_3_out, I0 =>  C_22_S_3_L_0_out, I1 =>  C_22_S_3_L_1_out, I2 =>  C_22_S_3_L_2_out, I3 =>  C_22_S_3_L_3_out, I4 =>  C_22_S_3_L_4_out, I5 =>  C_22_S_3_L_5_out); 
C_22_S_4_inst : LUT6 generic map(INIT => "1111111011111110111010001000100011101110111010001000000010000000") port map( O =>C_22_S_4_out, I0 =>  C_22_S_4_L_0_out, I1 =>  C_22_S_4_L_1_out, I2 =>  C_22_S_4_L_2_out, I3 =>  C_22_S_4_L_3_out, I4 =>  C_22_S_4_L_4_out, I5 =>  C_22_S_4_L_5_out); 
C_22_S_5_inst : LUT6 generic map(INIT => "1111111111101010111111101000000011111110100000001010100000000000") port map( O =>C_22_S_5_out, I0 =>  C_22_S_5_L_0_out, I1 =>  C_22_S_5_L_1_out, I2 =>  C_22_S_5_L_2_out, I3 =>  C_22_S_5_L_3_out, I4 =>  C_22_S_5_L_4_out, I5 =>  C_22_S_5_L_5_out); 

C_22_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_22_out, I0 =>  C_22_S_0_out, I1 =>  C_22_S_1_out, I2 =>  C_22_S_2_out, I3 =>  C_22_S_3_out, I4 =>  C_22_S_4_out, I5 =>  C_22_S_5_out); 

 
C_23_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_23_S_0_out, I0 =>  C_23_S_0_L_0_out, I1 =>  C_23_S_0_L_1_out, I2 =>  C_23_S_0_L_2_out, I3 =>  C_23_S_0_L_3_out, I4 =>  C_23_S_0_L_4_out, I5 =>  C_23_S_0_L_5_out); 
C_23_S_1_inst : LUT6 generic map(INIT => "1110111011101010111011101010100011101010100010001010100010001000") port map( O =>C_23_S_1_out, I0 =>  C_23_S_1_L_0_out, I1 =>  C_23_S_1_L_1_out, I2 =>  C_23_S_1_L_2_out, I3 =>  C_23_S_1_L_3_out, I4 =>  C_23_S_1_L_4_out, I5 =>  C_23_S_1_L_5_out); 
C_23_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_23_S_2_out, I0 =>  C_23_S_2_L_0_out, I1 =>  C_23_S_2_L_1_out, I2 =>  C_23_S_2_L_2_out, I3 =>  C_23_S_2_L_3_out, I4 =>  C_23_S_2_L_4_out, I5 =>  C_23_S_2_L_5_out); 
C_23_S_3_inst : LUT6 generic map(INIT => "1111111011111000111110001110000011111000111000001110000010000000") port map( O =>C_23_S_3_out, I0 =>  C_23_S_3_L_0_out, I1 =>  C_23_S_3_L_1_out, I2 =>  C_23_S_3_L_2_out, I3 =>  C_23_S_3_L_3_out, I4 =>  C_23_S_3_L_4_out, I5 =>  C_23_S_3_L_5_out); 
C_23_S_4_inst : LUT6 generic map(INIT => "1111111111101110111111101010100011101010100000001000100000000000") port map( O =>C_23_S_4_out, I0 =>  C_23_S_4_L_0_out, I1 =>  C_23_S_4_L_1_out, I2 =>  C_23_S_4_L_2_out, I3 =>  C_23_S_4_L_3_out, I4 =>  C_23_S_4_L_4_out, I5 =>  C_23_S_4_L_5_out); 
C_23_S_5_inst : LUT6 generic map(INIT => "1111111011101110111010101000100011101110101010001000100010000000") port map( O =>C_23_S_5_out, I0 =>  C_23_S_5_L_0_out, I1 =>  C_23_S_5_L_1_out, I2 =>  C_23_S_5_L_2_out, I3 =>  C_23_S_5_L_3_out, I4 =>  C_23_S_5_L_4_out, I5 =>  C_23_S_5_L_5_out); 

C_23_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_23_out, I0 =>  C_23_S_0_out, I1 =>  C_23_S_1_out, I2 =>  C_23_S_2_out, I3 =>  C_23_S_3_out, I4 =>  C_23_S_4_out, I5 =>  C_23_S_5_out); 

 
C_24_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_24_S_0_out, I0 =>  C_24_S_0_L_0_out, I1 =>  C_24_S_0_L_1_out, I2 =>  C_24_S_0_L_2_out, I3 =>  C_24_S_0_L_3_out, I4 =>  C_24_S_0_L_4_out, I5 =>  C_24_S_0_L_5_out); 
C_24_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_24_S_1_out, I0 =>  C_24_S_1_L_0_out, I1 =>  C_24_S_1_L_1_out, I2 =>  C_24_S_1_L_2_out, I3 =>  C_24_S_1_L_3_out, I4 =>  C_24_S_1_L_4_out, I5 =>  C_24_S_1_L_5_out); 
C_24_S_2_inst : LUT6 generic map(INIT => "1111111011101010111111101010100011101010100000001010100010000000") port map( O =>C_24_S_2_out, I0 =>  C_24_S_2_L_0_out, I1 =>  C_24_S_2_L_1_out, I2 =>  C_24_S_2_L_2_out, I3 =>  C_24_S_2_L_3_out, I4 =>  C_24_S_2_L_4_out, I5 =>  C_24_S_2_L_5_out); 
C_24_S_3_inst : LUT6 generic map(INIT => "1111111111111110111011001100100011101100110010001000000000000000") port map( O =>C_24_S_3_out, I0 =>  C_24_S_3_L_0_out, I1 =>  C_24_S_3_L_1_out, I2 =>  C_24_S_3_L_2_out, I3 =>  C_24_S_3_L_3_out, I4 =>  C_24_S_3_L_4_out, I5 =>  C_24_S_3_L_5_out); 
C_24_S_4_inst : LUT6 generic map(INIT => "1111111011101100111011101100100011101100100010001100100010000000") port map( O =>C_24_S_4_out, I0 =>  C_24_S_4_L_0_out, I1 =>  C_24_S_4_L_1_out, I2 =>  C_24_S_4_L_2_out, I3 =>  C_24_S_4_L_3_out, I4 =>  C_24_S_4_L_4_out, I5 =>  C_24_S_4_L_5_out); 
C_24_S_5_inst : LUT6 generic map(INIT => "1111111011101110111011101110100011101000100010001000100010000000") port map( O =>C_24_S_5_out, I0 =>  C_24_S_5_L_0_out, I1 =>  C_24_S_5_L_1_out, I2 =>  C_24_S_5_L_2_out, I3 =>  C_24_S_5_L_3_out, I4 =>  C_24_S_5_L_4_out, I5 =>  C_24_S_5_L_5_out); 

C_24_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_24_out, I0 =>  C_24_S_0_out, I1 =>  C_24_S_1_out, I2 =>  C_24_S_2_out, I3 =>  C_24_S_3_out, I4 =>  C_24_S_4_out, I5 =>  C_24_S_5_out); 

 
C_25_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_25_S_0_out, I0 =>  C_25_S_0_L_0_out, I1 =>  C_25_S_0_L_1_out, I2 =>  C_25_S_0_L_2_out, I3 =>  C_25_S_0_L_3_out, I4 =>  C_25_S_0_L_4_out, I5 =>  C_25_S_0_L_5_out); 
C_25_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101110100011101000101010001010100010000000") port map( O =>C_25_S_1_out, I0 =>  C_25_S_1_L_0_out, I1 =>  C_25_S_1_L_1_out, I2 =>  C_25_S_1_L_2_out, I3 =>  C_25_S_1_L_3_out, I4 =>  C_25_S_1_L_4_out, I5 =>  C_25_S_1_L_5_out); 
C_25_S_2_inst : LUT6 generic map(INIT => "1111111111111110111111101010100011101010100000001000000000000000") port map( O =>C_25_S_2_out, I0 =>  C_25_S_2_L_0_out, I1 =>  C_25_S_2_L_1_out, I2 =>  C_25_S_2_L_2_out, I3 =>  C_25_S_2_L_3_out, I4 =>  C_25_S_2_L_4_out, I5 =>  C_25_S_2_L_5_out); 
C_25_S_3_inst : LUT6 generic map(INIT => "1111111111111110111010001000000011111110111010001000000000000000") port map( O =>C_25_S_3_out, I0 =>  C_25_S_3_L_0_out, I1 =>  C_25_S_3_L_1_out, I2 =>  C_25_S_3_L_2_out, I3 =>  C_25_S_3_L_3_out, I4 =>  C_25_S_3_L_4_out, I5 =>  C_25_S_3_L_5_out); 
C_25_S_4_inst : LUT6 generic map(INIT => "1111111111111110111011001100000011111100110010001000000000000000") port map( O =>C_25_S_4_out, I0 =>  C_25_S_4_L_0_out, I1 =>  C_25_S_4_L_1_out, I2 =>  C_25_S_4_L_2_out, I3 =>  C_25_S_4_L_3_out, I4 =>  C_25_S_4_L_4_out, I5 =>  C_25_S_4_L_5_out); 
C_25_S_5_inst : LUT6 generic map(INIT => "1111111111101100111111101100000011111100100000001100100000000000") port map( O =>C_25_S_5_out, I0 =>  C_25_S_5_L_0_out, I1 =>  C_25_S_5_L_1_out, I2 =>  C_25_S_5_L_2_out, I3 =>  C_25_S_5_L_3_out, I4 =>  C_25_S_5_L_4_out, I5 =>  C_25_S_5_L_5_out); 

C_25_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_25_out, I0 =>  C_25_S_0_out, I1 =>  C_25_S_1_out, I2 =>  C_25_S_2_out, I3 =>  C_25_S_3_out, I4 =>  C_25_S_4_out, I5 =>  C_25_S_5_out); 

 
C_26_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_26_S_0_out, I0 =>  C_26_S_0_L_0_out, I1 =>  C_26_S_0_L_1_out, I2 =>  C_26_S_0_L_2_out, I3 =>  C_26_S_0_L_3_out, I4 =>  C_26_S_0_L_4_out, I5 =>  C_26_S_0_L_5_out); 
C_26_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_26_S_1_out, I0 =>  C_26_S_1_L_0_out, I1 =>  C_26_S_1_L_1_out, I2 =>  C_26_S_1_L_2_out, I3 =>  C_26_S_1_L_3_out, I4 =>  C_26_S_1_L_4_out, I5 =>  C_26_S_1_L_5_out); 
C_26_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_26_S_2_out, I0 =>  C_26_S_2_L_0_out, I1 =>  C_26_S_2_L_1_out, I2 =>  C_26_S_2_L_2_out, I3 =>  C_26_S_2_L_3_out, I4 =>  C_26_S_2_L_4_out, I5 =>  C_26_S_2_L_5_out); 
C_26_S_3_inst : LUT6 generic map(INIT => "1111111111111100111111001110000011111000110000001100000000000000") port map( O =>C_26_S_3_out, I0 =>  C_26_S_3_L_0_out, I1 =>  C_26_S_3_L_1_out, I2 =>  C_26_S_3_L_2_out, I3 =>  C_26_S_3_L_3_out, I4 =>  C_26_S_3_L_4_out, I5 =>  C_26_S_3_L_5_out); 
C_26_S_4_inst : LUT6 generic map(INIT => "1111111111111010111111101010100011101010100000001010000000000000") port map( O =>C_26_S_4_out, I0 =>  C_26_S_4_L_0_out, I1 =>  C_26_S_4_L_1_out, I2 =>  C_26_S_4_L_2_out, I3 =>  C_26_S_4_L_3_out, I4 =>  C_26_S_4_L_4_out, I5 =>  C_26_S_4_L_5_out); 
C_26_S_5_inst : LUT6 generic map(INIT => "1111111011111010111110101110100011101000101000001010000010000000") port map( O =>C_26_S_5_out, I0 =>  C_26_S_5_L_0_out, I1 =>  C_26_S_5_L_1_out, I2 =>  C_26_S_5_L_2_out, I3 =>  C_26_S_5_L_3_out, I4 =>  C_26_S_5_L_4_out, I5 =>  C_26_S_5_L_5_out); 

C_26_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_26_out, I0 =>  C_26_S_0_out, I1 =>  C_26_S_1_out, I2 =>  C_26_S_2_out, I3 =>  C_26_S_3_out, I4 =>  C_26_S_4_out, I5 =>  C_26_S_5_out); 

 
C_27_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_27_S_0_out, I0 =>  C_27_S_0_L_0_out, I1 =>  C_27_S_0_L_1_out, I2 =>  C_27_S_0_L_2_out, I3 =>  C_27_S_0_L_3_out, I4 =>  C_27_S_0_L_4_out, I5 =>  C_27_S_0_L_5_out); 
C_27_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101110100011101000101010001010100010000000") port map( O =>C_27_S_1_out, I0 =>  C_27_S_1_L_0_out, I1 =>  C_27_S_1_L_1_out, I2 =>  C_27_S_1_L_2_out, I3 =>  C_27_S_1_L_3_out, I4 =>  C_27_S_1_L_4_out, I5 =>  C_27_S_1_L_5_out); 
C_27_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001110100011101000111010001110100010000000") port map( O =>C_27_S_2_out, I0 =>  C_27_S_2_L_0_out, I1 =>  C_27_S_2_L_1_out, I2 =>  C_27_S_2_L_2_out, I3 =>  C_27_S_2_L_3_out, I4 =>  C_27_S_2_L_4_out, I5 =>  C_27_S_2_L_5_out); 
C_27_S_3_inst : LUT6 generic map(INIT => "1111111011111110111010001100100011101100111010001000000010000000") port map( O =>C_27_S_3_out, I0 =>  C_27_S_3_L_0_out, I1 =>  C_27_S_3_L_1_out, I2 =>  C_27_S_3_L_2_out, I3 =>  C_27_S_3_L_3_out, I4 =>  C_27_S_3_L_4_out, I5 =>  C_27_S_3_L_5_out); 
C_27_S_4_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_27_S_4_out, I0 =>  C_27_S_4_L_0_out, I1 =>  C_27_S_4_L_1_out, I2 =>  C_27_S_4_L_2_out, I3 =>  C_27_S_4_L_3_out, I4 =>  C_27_S_4_L_4_out, I5 =>  C_27_S_4_L_5_out); 
C_27_S_5_inst : LUT6 generic map(INIT => "1111111011101000111011101000000011111110100010001110100010000000") port map( O =>C_27_S_5_out, I0 =>  C_27_S_5_L_0_out, I1 =>  C_27_S_5_L_1_out, I2 =>  C_27_S_5_L_2_out, I3 =>  C_27_S_5_L_3_out, I4 =>  C_27_S_5_L_4_out, I5 =>  C_27_S_5_L_5_out); 

C_27_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_27_out, I0 =>  C_27_S_0_out, I1 =>  C_27_S_1_out, I2 =>  C_27_S_2_out, I3 =>  C_27_S_3_out, I4 =>  C_27_S_4_out, I5 =>  C_27_S_5_out); 

 
C_28_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_28_S_0_out, I0 =>  C_28_S_0_L_0_out, I1 =>  C_28_S_0_L_1_out, I2 =>  C_28_S_0_L_2_out, I3 =>  C_28_S_0_L_3_out, I4 =>  C_28_S_0_L_4_out, I5 =>  C_28_S_0_L_5_out); 
C_28_S_1_inst : LUT6 generic map(INIT => "1110101011101010101010101010100011101010101010101010100010101000") port map( O =>C_28_S_1_out, I0 =>  C_28_S_1_L_0_out, I1 =>  C_28_S_1_L_1_out, I2 =>  C_28_S_1_L_2_out, I3 =>  C_28_S_1_L_3_out, I4 =>  C_28_S_1_L_4_out, I5 =>  C_28_S_1_L_5_out); 
C_28_S_2_inst : LUT6 generic map(INIT => "1111111011111100111111001110100011101000110000001100000010000000") port map( O =>C_28_S_2_out, I0 =>  C_28_S_2_L_0_out, I1 =>  C_28_S_2_L_1_out, I2 =>  C_28_S_2_L_2_out, I3 =>  C_28_S_2_L_3_out, I4 =>  C_28_S_2_L_4_out, I5 =>  C_28_S_2_L_5_out); 
C_28_S_3_inst : LUT6 generic map(INIT => "1111111111101010111010101000000011111110101010001010100000000000") port map( O =>C_28_S_3_out, I0 =>  C_28_S_3_L_0_out, I1 =>  C_28_S_3_L_1_out, I2 =>  C_28_S_3_L_2_out, I3 =>  C_28_S_3_L_3_out, I4 =>  C_28_S_3_L_4_out, I5 =>  C_28_S_3_L_5_out); 
C_28_S_4_inst : LUT6 generic map(INIT => "1111111111101000111111101110100011101000100000001110100000000000") port map( O =>C_28_S_4_out, I0 =>  C_28_S_4_L_0_out, I1 =>  C_28_S_4_L_1_out, I2 =>  C_28_S_4_L_2_out, I3 =>  C_28_S_4_L_3_out, I4 =>  C_28_S_4_L_4_out, I5 =>  C_28_S_4_L_5_out); 
C_28_S_5_inst : LUT6 generic map(INIT => "1111111111101010111110101010100011101010101000001010100000000000") port map( O =>C_28_S_5_out, I0 =>  C_28_S_5_L_0_out, I1 =>  C_28_S_5_L_1_out, I2 =>  C_28_S_5_L_2_out, I3 =>  C_28_S_5_L_3_out, I4 =>  C_28_S_5_L_4_out, I5 =>  C_28_S_5_L_5_out); 

C_28_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_28_out, I0 =>  C_28_S_0_out, I1 =>  C_28_S_1_out, I2 =>  C_28_S_2_out, I3 =>  C_28_S_3_out, I4 =>  C_28_S_4_out, I5 =>  C_28_S_5_out); 

 
C_29_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_29_S_0_out, I0 =>  C_29_S_0_L_0_out, I1 =>  C_29_S_0_L_1_out, I2 =>  C_29_S_0_L_2_out, I3 =>  C_29_S_0_L_3_out, I4 =>  C_29_S_0_L_4_out, I5 =>  C_29_S_0_L_5_out); 
C_29_S_1_inst : LUT6 generic map(INIT => "1110111011101000111011001100100011101100110010001110100010001000") port map( O =>C_29_S_1_out, I0 =>  C_29_S_1_L_0_out, I1 =>  C_29_S_1_L_1_out, I2 =>  C_29_S_1_L_2_out, I3 =>  C_29_S_1_L_3_out, I4 =>  C_29_S_1_L_4_out, I5 =>  C_29_S_1_L_5_out); 
C_29_S_2_inst : LUT6 generic map(INIT => "1111111011101000111111101100100011101100100000001110100010000000") port map( O =>C_29_S_2_out, I0 =>  C_29_S_2_L_0_out, I1 =>  C_29_S_2_L_1_out, I2 =>  C_29_S_2_L_2_out, I3 =>  C_29_S_2_L_3_out, I4 =>  C_29_S_2_L_4_out, I5 =>  C_29_S_2_L_5_out); 
C_29_S_3_inst : LUT6 generic map(INIT => "1111111111101010111111101010100011101010100000001010100000000000") port map( O =>C_29_S_3_out, I0 =>  C_29_S_3_L_0_out, I1 =>  C_29_S_3_L_1_out, I2 =>  C_29_S_3_L_2_out, I3 =>  C_29_S_3_L_3_out, I4 =>  C_29_S_3_L_4_out, I5 =>  C_29_S_3_L_5_out); 
C_29_S_4_inst : LUT6 generic map(INIT => "1111111011101110111011101100100011101100100010001000100010000000") port map( O =>C_29_S_4_out, I0 =>  C_29_S_4_L_0_out, I1 =>  C_29_S_4_L_1_out, I2 =>  C_29_S_4_L_2_out, I3 =>  C_29_S_4_L_3_out, I4 =>  C_29_S_4_L_4_out, I5 =>  C_29_S_4_L_5_out); 
C_29_S_5_inst : LUT6 generic map(INIT => "1111111011101010111110101010000011111010101000001010100010000000") port map( O =>C_29_S_5_out, I0 =>  C_29_S_5_L_0_out, I1 =>  C_29_S_5_L_1_out, I2 =>  C_29_S_5_L_2_out, I3 =>  C_29_S_5_L_3_out, I4 =>  C_29_S_5_L_4_out, I5 =>  C_29_S_5_L_5_out); 

C_29_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_29_out, I0 =>  C_29_S_0_out, I1 =>  C_29_S_1_out, I2 =>  C_29_S_2_out, I3 =>  C_29_S_3_out, I4 =>  C_29_S_4_out, I5 =>  C_29_S_5_out); 

 
C_30_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_30_S_0_out, I0 =>  C_30_S_0_L_0_out, I1 =>  C_30_S_0_L_1_out, I2 =>  C_30_S_0_L_2_out, I3 =>  C_30_S_0_L_3_out, I4 =>  C_30_S_0_L_4_out, I5 =>  C_30_S_0_L_5_out); 
C_30_S_1_inst : LUT6 generic map(INIT => "1111101011101010111010101010100011101010101010001010100010100000") port map( O =>C_30_S_1_out, I0 =>  C_30_S_1_L_0_out, I1 =>  C_30_S_1_L_1_out, I2 =>  C_30_S_1_L_2_out, I3 =>  C_30_S_1_L_3_out, I4 =>  C_30_S_1_L_4_out, I5 =>  C_30_S_1_L_5_out); 
C_30_S_2_inst : LUT6 generic map(INIT => "1111111011111000111110101010000011111010101000001110000010000000") port map( O =>C_30_S_2_out, I0 =>  C_30_S_2_L_0_out, I1 =>  C_30_S_2_L_1_out, I2 =>  C_30_S_2_L_2_out, I3 =>  C_30_S_2_L_3_out, I4 =>  C_30_S_2_L_4_out, I5 =>  C_30_S_2_L_5_out); 
C_30_S_3_inst : LUT6 generic map(INIT => "1111111111101100111011101000100011101110100010001100100000000000") port map( O =>C_30_S_3_out, I0 =>  C_30_S_3_L_0_out, I1 =>  C_30_S_3_L_1_out, I2 =>  C_30_S_3_L_2_out, I3 =>  C_30_S_3_L_3_out, I4 =>  C_30_S_3_L_4_out, I5 =>  C_30_S_3_L_5_out); 
C_30_S_4_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_30_S_4_out, I0 =>  C_30_S_4_L_0_out, I1 =>  C_30_S_4_L_1_out, I2 =>  C_30_S_4_L_2_out, I3 =>  C_30_S_4_L_3_out, I4 =>  C_30_S_4_L_4_out, I5 =>  C_30_S_4_L_5_out); 
C_30_S_5_inst : LUT6 generic map(INIT => "1111111111101110111011001100100011101100110010001000100000000000") port map( O =>C_30_S_5_out, I0 =>  C_30_S_5_L_0_out, I1 =>  C_30_S_5_L_1_out, I2 =>  C_30_S_5_L_2_out, I3 =>  C_30_S_5_L_3_out, I4 =>  C_30_S_5_L_4_out, I5 =>  C_30_S_5_L_5_out); 

C_30_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_30_out, I0 =>  C_30_S_0_out, I1 =>  C_30_S_1_out, I2 =>  C_30_S_2_out, I3 =>  C_30_S_3_out, I4 =>  C_30_S_4_out, I5 =>  C_30_S_5_out); 

 
C_31_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_31_S_0_out, I0 =>  C_31_S_0_L_0_out, I1 =>  C_31_S_0_L_1_out, I2 =>  C_31_S_0_L_2_out, I3 =>  C_31_S_0_L_3_out, I4 =>  C_31_S_0_L_4_out, I5 =>  C_31_S_0_L_5_out); 
C_31_S_1_inst : LUT6 generic map(INIT => "1110101011101010111010001010100011101010111010001010100010101000") port map( O =>C_31_S_1_out, I0 =>  C_31_S_1_L_0_out, I1 =>  C_31_S_1_L_1_out, I2 =>  C_31_S_1_L_2_out, I3 =>  C_31_S_1_L_3_out, I4 =>  C_31_S_1_L_4_out, I5 =>  C_31_S_1_L_5_out); 
C_31_S_2_inst : LUT6 generic map(INIT => "1111111011101000111011101000100011101110100010001110100010000000") port map( O =>C_31_S_2_out, I0 =>  C_31_S_2_L_0_out, I1 =>  C_31_S_2_L_1_out, I2 =>  C_31_S_2_L_2_out, I3 =>  C_31_S_2_L_3_out, I4 =>  C_31_S_2_L_4_out, I5 =>  C_31_S_2_L_5_out); 
C_31_S_3_inst : LUT6 generic map(INIT => "1111111111111110111010001000000011111110111010001000000000000000") port map( O =>C_31_S_3_out, I0 =>  C_31_S_3_L_0_out, I1 =>  C_31_S_3_L_1_out, I2 =>  C_31_S_3_L_2_out, I3 =>  C_31_S_3_L_3_out, I4 =>  C_31_S_3_L_4_out, I5 =>  C_31_S_3_L_5_out); 
C_31_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010101000100011101110101010001010100010000000") port map( O =>C_31_S_4_out, I0 =>  C_31_S_4_L_0_out, I1 =>  C_31_S_4_L_1_out, I2 =>  C_31_S_4_L_2_out, I3 =>  C_31_S_4_L_3_out, I4 =>  C_31_S_4_L_4_out, I5 =>  C_31_S_4_L_5_out); 
C_31_S_5_inst : LUT6 generic map(INIT => "1111111111111000111110001000000011111110111000001110000000000000") port map( O =>C_31_S_5_out, I0 =>  C_31_S_5_L_0_out, I1 =>  C_31_S_5_L_1_out, I2 =>  C_31_S_5_L_2_out, I3 =>  C_31_S_5_L_3_out, I4 =>  C_31_S_5_L_4_out, I5 =>  C_31_S_5_L_5_out); 

C_31_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_31_out, I0 =>  C_31_S_0_out, I1 =>  C_31_S_1_out, I2 =>  C_31_S_2_out, I3 =>  C_31_S_3_out, I4 =>  C_31_S_4_out, I5 =>  C_31_S_5_out); 

 
C_32_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_32_S_0_out, I0 =>  C_32_S_0_L_0_out, I1 =>  C_32_S_0_L_1_out, I2 =>  C_32_S_0_L_2_out, I3 =>  C_32_S_0_L_3_out, I4 =>  C_32_S_0_L_4_out, I5 =>  C_32_S_0_L_5_out); 
C_32_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_32_S_1_out, I0 =>  C_32_S_1_L_0_out, I1 =>  C_32_S_1_L_1_out, I2 =>  C_32_S_1_L_2_out, I3 =>  C_32_S_1_L_3_out, I4 =>  C_32_S_1_L_4_out, I5 =>  C_32_S_1_L_5_out); 
C_32_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010001010100011101010111010001010100010000000") port map( O =>C_32_S_2_out, I0 =>  C_32_S_2_L_0_out, I1 =>  C_32_S_2_L_1_out, I2 =>  C_32_S_2_L_2_out, I3 =>  C_32_S_2_L_3_out, I4 =>  C_32_S_2_L_4_out, I5 =>  C_32_S_2_L_5_out); 
C_32_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001010100011101010111010001110100010000000") port map( O =>C_32_S_3_out, I0 =>  C_32_S_3_L_0_out, I1 =>  C_32_S_3_L_1_out, I2 =>  C_32_S_3_L_2_out, I3 =>  C_32_S_3_L_3_out, I4 =>  C_32_S_3_L_4_out, I5 =>  C_32_S_3_L_5_out); 
C_32_S_4_inst : LUT6 generic map(INIT => "1111111011101000111011101000100011101110100010001110100010000000") port map( O =>C_32_S_4_out, I0 =>  C_32_S_4_L_0_out, I1 =>  C_32_S_4_L_1_out, I2 =>  C_32_S_4_L_2_out, I3 =>  C_32_S_4_L_3_out, I4 =>  C_32_S_4_L_4_out, I5 =>  C_32_S_4_L_5_out); 
C_32_S_5_inst : LUT6 generic map(INIT => "1111111011101000111011101000100011101110100010001110100010000000") port map( O =>C_32_S_5_out, I0 =>  C_32_S_5_L_0_out, I1 =>  C_32_S_5_L_1_out, I2 =>  C_32_S_5_L_2_out, I3 =>  C_32_S_5_L_3_out, I4 =>  C_32_S_5_L_4_out, I5 =>  C_32_S_5_L_5_out); 

C_32_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_32_out, I0 =>  C_32_S_0_out, I1 =>  C_32_S_1_out, I2 =>  C_32_S_2_out, I3 =>  C_32_S_3_out, I4 =>  C_32_S_4_out, I5 =>  C_32_S_5_out); 

 
C_33_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_33_S_0_out, I0 =>  C_33_S_0_L_0_out, I1 =>  C_33_S_0_L_1_out, I2 =>  C_33_S_0_L_2_out, I3 =>  C_33_S_0_L_3_out, I4 =>  C_33_S_0_L_4_out, I5 =>  C_33_S_0_L_5_out); 
C_33_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_33_S_1_out, I0 =>  C_33_S_1_L_0_out, I1 =>  C_33_S_1_L_1_out, I2 =>  C_33_S_1_L_2_out, I3 =>  C_33_S_1_L_3_out, I4 =>  C_33_S_1_L_4_out, I5 =>  C_33_S_1_L_5_out); 
C_33_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010101010000011111010101010001110100010000000") port map( O =>C_33_S_2_out, I0 =>  C_33_S_2_L_0_out, I1 =>  C_33_S_2_L_1_out, I2 =>  C_33_S_2_L_2_out, I3 =>  C_33_S_2_L_3_out, I4 =>  C_33_S_2_L_4_out, I5 =>  C_33_S_2_L_5_out); 
C_33_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001110100011101000111010001110100010000000") port map( O =>C_33_S_3_out, I0 =>  C_33_S_3_L_0_out, I1 =>  C_33_S_3_L_1_out, I2 =>  C_33_S_3_L_2_out, I3 =>  C_33_S_3_L_3_out, I4 =>  C_33_S_3_L_4_out, I5 =>  C_33_S_3_L_5_out); 
C_33_S_4_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_33_S_4_out, I0 =>  C_33_S_4_L_0_out, I1 =>  C_33_S_4_L_1_out, I2 =>  C_33_S_4_L_2_out, I3 =>  C_33_S_4_L_3_out, I4 =>  C_33_S_4_L_4_out, I5 =>  C_33_S_4_L_5_out); 
C_33_S_5_inst : LUT6 generic map(INIT => "1111111011111000111010001010000011111010111010001110000010000000") port map( O =>C_33_S_5_out, I0 =>  C_33_S_5_L_0_out, I1 =>  C_33_S_5_L_1_out, I2 =>  C_33_S_5_L_2_out, I3 =>  C_33_S_5_L_3_out, I4 =>  C_33_S_5_L_4_out, I5 =>  C_33_S_5_L_5_out); 

C_33_inst : LUT6 generic map(INIT => "1110101010101010111010101010101010101010101010001010101010101000") port map( O =>C_33_out, I0 =>  C_33_S_0_out, I1 =>  C_33_S_1_out, I2 =>  C_33_S_2_out, I3 =>  C_33_S_3_out, I4 =>  C_33_S_4_out, I5 =>  C_33_S_5_out); 

 
C_34_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_34_S_0_out, I0 =>  C_34_S_0_L_0_out, I1 =>  C_34_S_0_L_1_out, I2 =>  C_34_S_0_L_2_out, I3 =>  C_34_S_0_L_3_out, I4 =>  C_34_S_0_L_4_out, I5 =>  C_34_S_0_L_5_out); 
C_34_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010001010100011101010111010001010100010000000") port map( O =>C_34_S_1_out, I0 =>  C_34_S_1_L_0_out, I1 =>  C_34_S_1_L_1_out, I2 =>  C_34_S_1_L_2_out, I3 =>  C_34_S_1_L_3_out, I4 =>  C_34_S_1_L_4_out, I5 =>  C_34_S_1_L_5_out); 
C_34_S_2_inst : LUT6 generic map(INIT => "1111111011111100111010001100000011111100111010001100000010000000") port map( O =>C_34_S_2_out, I0 =>  C_34_S_2_L_0_out, I1 =>  C_34_S_2_L_1_out, I2 =>  C_34_S_2_L_2_out, I3 =>  C_34_S_2_L_3_out, I4 =>  C_34_S_2_L_4_out, I5 =>  C_34_S_2_L_5_out); 
C_34_S_3_inst : LUT6 generic map(INIT => "1111111011111100111110001110100011101000111000001100000010000000") port map( O =>C_34_S_3_out, I0 =>  C_34_S_3_L_0_out, I1 =>  C_34_S_3_L_1_out, I2 =>  C_34_S_3_L_2_out, I3 =>  C_34_S_3_L_3_out, I4 =>  C_34_S_3_L_4_out, I5 =>  C_34_S_3_L_5_out); 
C_34_S_4_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_34_S_4_out, I0 =>  C_34_S_4_L_0_out, I1 =>  C_34_S_4_L_1_out, I2 =>  C_34_S_4_L_2_out, I3 =>  C_34_S_4_L_3_out, I4 =>  C_34_S_4_L_4_out, I5 =>  C_34_S_4_L_5_out); 
C_34_S_5_inst : LUT6 generic map(INIT => "1111111011101000111110101010000011111010101000001110100010000000") port map( O =>C_34_S_5_out, I0 =>  C_34_S_5_L_0_out, I1 =>  C_34_S_5_L_1_out, I2 =>  C_34_S_5_L_2_out, I3 =>  C_34_S_5_L_3_out, I4 =>  C_34_S_5_L_4_out, I5 =>  C_34_S_5_L_5_out); 

C_34_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_34_out, I0 =>  C_34_S_0_out, I1 =>  C_34_S_1_out, I2 =>  C_34_S_2_out, I3 =>  C_34_S_3_out, I4 =>  C_34_S_4_out, I5 =>  C_34_S_5_out); 

 
C_35_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_35_S_0_out, I0 =>  C_35_S_0_L_0_out, I1 =>  C_35_S_0_L_1_out, I2 =>  C_35_S_0_L_2_out, I3 =>  C_35_S_0_L_3_out, I4 =>  C_35_S_0_L_4_out, I5 =>  C_35_S_0_L_5_out); 
C_35_S_1_inst : LUT6 generic map(INIT => "1111111010101010111010101010100011101010101010001010101010000000") port map( O =>C_35_S_1_out, I0 =>  C_35_S_1_L_0_out, I1 =>  C_35_S_1_L_1_out, I2 =>  C_35_S_1_L_2_out, I3 =>  C_35_S_1_L_3_out, I4 =>  C_35_S_1_L_4_out, I5 =>  C_35_S_1_L_5_out); 
C_35_S_2_inst : LUT6 generic map(INIT => "1111111011111000111110001110000011111000111000001110000010000000") port map( O =>C_35_S_2_out, I0 =>  C_35_S_2_L_0_out, I1 =>  C_35_S_2_L_1_out, I2 =>  C_35_S_2_L_2_out, I3 =>  C_35_S_2_L_3_out, I4 =>  C_35_S_2_L_4_out, I5 =>  C_35_S_2_L_5_out); 
C_35_S_3_inst : LUT6 generic map(INIT => "1111111011101010111010001010100011101010111010001010100010000000") port map( O =>C_35_S_3_out, I0 =>  C_35_S_3_L_0_out, I1 =>  C_35_S_3_L_1_out, I2 =>  C_35_S_3_L_2_out, I3 =>  C_35_S_3_L_3_out, I4 =>  C_35_S_3_L_4_out, I5 =>  C_35_S_3_L_5_out); 
C_35_S_4_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_35_S_4_out, I0 =>  C_35_S_4_L_0_out, I1 =>  C_35_S_4_L_1_out, I2 =>  C_35_S_4_L_2_out, I3 =>  C_35_S_4_L_3_out, I4 =>  C_35_S_4_L_4_out, I5 =>  C_35_S_4_L_5_out); 
C_35_S_5_inst : LUT6 generic map(INIT => "1111111111101100111011001000000011111110110010001100100000000000") port map( O =>C_35_S_5_out, I0 =>  C_35_S_5_L_0_out, I1 =>  C_35_S_5_L_1_out, I2 =>  C_35_S_5_L_2_out, I3 =>  C_35_S_5_L_3_out, I4 =>  C_35_S_5_L_4_out, I5 =>  C_35_S_5_L_5_out); 

C_35_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_35_out, I0 =>  C_35_S_0_out, I1 =>  C_35_S_1_out, I2 =>  C_35_S_2_out, I3 =>  C_35_S_3_out, I4 =>  C_35_S_4_out, I5 =>  C_35_S_5_out); 

 
C_36_S_0_inst : LUT6 generic map(INIT => "1110111011101010101010101010100011101010101010101010100010001000") port map( O =>C_36_S_0_out, I0 =>  C_36_S_0_L_0_out, I1 =>  C_36_S_0_L_1_out, I2 =>  C_36_S_0_L_2_out, I3 =>  C_36_S_0_L_3_out, I4 =>  C_36_S_0_L_4_out, I5 =>  C_36_S_0_L_5_out); 
C_36_S_1_inst : LUT6 generic map(INIT => "1111111111101110111011101010100011101010100010001000100000000000") port map( O =>C_36_S_1_out, I0 =>  C_36_S_1_L_0_out, I1 =>  C_36_S_1_L_1_out, I2 =>  C_36_S_1_L_2_out, I3 =>  C_36_S_1_L_3_out, I4 =>  C_36_S_1_L_4_out, I5 =>  C_36_S_1_L_5_out); 
C_36_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101000100011101110101010001010100010000000") port map( O =>C_36_S_2_out, I0 =>  C_36_S_2_L_0_out, I1 =>  C_36_S_2_L_1_out, I2 =>  C_36_S_2_L_2_out, I3 =>  C_36_S_2_L_3_out, I4 =>  C_36_S_2_L_4_out, I5 =>  C_36_S_2_L_5_out); 
C_36_S_3_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_36_S_3_out, I0 =>  C_36_S_3_L_0_out, I1 =>  C_36_S_3_L_1_out, I2 =>  C_36_S_3_L_2_out, I3 =>  C_36_S_3_L_3_out, I4 =>  C_36_S_3_L_4_out, I5 =>  C_36_S_3_L_5_out); 
C_36_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_36_S_4_out, I0 =>  C_36_S_4_L_0_out, I1 =>  C_36_S_4_L_1_out, I2 =>  C_36_S_4_L_2_out, I3 =>  C_36_S_4_L_3_out, I4 =>  C_36_S_4_L_4_out, I5 =>  C_36_S_4_L_5_out); 
C_36_S_5_inst : LUT6 generic map(INIT => "1111111111111110111110001000000011111110111000001000000000000000") port map( O =>C_36_S_5_out, I0 =>  C_36_S_5_L_0_out, I1 =>  C_36_S_5_L_1_out, I2 =>  C_36_S_5_L_2_out, I3 =>  C_36_S_5_L_3_out, I4 =>  C_36_S_5_L_4_out, I5 =>  C_36_S_5_L_5_out); 

C_36_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_36_out, I0 =>  C_36_S_0_out, I1 =>  C_36_S_1_out, I2 =>  C_36_S_2_out, I3 =>  C_36_S_3_out, I4 =>  C_36_S_4_out, I5 =>  C_36_S_5_out); 

 
C_37_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_37_S_0_out, I0 =>  C_37_S_0_L_0_out, I1 =>  C_37_S_0_L_1_out, I2 =>  C_37_S_0_L_2_out, I3 =>  C_37_S_0_L_3_out, I4 =>  C_37_S_0_L_4_out, I5 =>  C_37_S_0_L_5_out); 
C_37_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010001110100011101000111010001010100010000000") port map( O =>C_37_S_1_out, I0 =>  C_37_S_1_L_0_out, I1 =>  C_37_S_1_L_1_out, I2 =>  C_37_S_1_L_2_out, I3 =>  C_37_S_1_L_3_out, I4 =>  C_37_S_1_L_4_out, I5 =>  C_37_S_1_L_5_out); 
C_37_S_2_inst : LUT6 generic map(INIT => "1111111011101110111010001000100011101110111010001000100010000000") port map( O =>C_37_S_2_out, I0 =>  C_37_S_2_L_0_out, I1 =>  C_37_S_2_L_1_out, I2 =>  C_37_S_2_L_2_out, I3 =>  C_37_S_2_L_3_out, I4 =>  C_37_S_2_L_4_out, I5 =>  C_37_S_2_L_5_out); 
C_37_S_3_inst : LUT6 generic map(INIT => "1111111111111110111011001100100011101100110010001000000000000000") port map( O =>C_37_S_3_out, I0 =>  C_37_S_3_L_0_out, I1 =>  C_37_S_3_L_1_out, I2 =>  C_37_S_3_L_2_out, I3 =>  C_37_S_3_L_3_out, I4 =>  C_37_S_3_L_4_out, I5 =>  C_37_S_3_L_5_out); 
C_37_S_4_inst : LUT6 generic map(INIT => "1111111011101000111111101110000011111000100000001110100010000000") port map( O =>C_37_S_4_out, I0 =>  C_37_S_4_L_0_out, I1 =>  C_37_S_4_L_1_out, I2 =>  C_37_S_4_L_2_out, I3 =>  C_37_S_4_L_3_out, I4 =>  C_37_S_4_L_4_out, I5 =>  C_37_S_4_L_5_out); 
C_37_S_5_inst : LUT6 generic map(INIT => "1111111111111010111010101010000011111010101010001010000000000000") port map( O =>C_37_S_5_out, I0 =>  C_37_S_5_L_0_out, I1 =>  C_37_S_5_L_1_out, I2 =>  C_37_S_5_L_2_out, I3 =>  C_37_S_5_L_3_out, I4 =>  C_37_S_5_L_4_out, I5 =>  C_37_S_5_L_5_out); 

C_37_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_37_out, I0 =>  C_37_S_0_out, I1 =>  C_37_S_1_out, I2 =>  C_37_S_2_out, I3 =>  C_37_S_3_out, I4 =>  C_37_S_4_out, I5 =>  C_37_S_5_out); 

 
C_38_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_38_S_0_out, I0 =>  C_38_S_0_L_0_out, I1 =>  C_38_S_0_L_1_out, I2 =>  C_38_S_0_L_2_out, I3 =>  C_38_S_0_L_3_out, I4 =>  C_38_S_0_L_4_out, I5 =>  C_38_S_0_L_5_out); 
C_38_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010001110100011101000111010001110100010000000") port map( O =>C_38_S_1_out, I0 =>  C_38_S_1_L_0_out, I1 =>  C_38_S_1_L_1_out, I2 =>  C_38_S_1_L_2_out, I3 =>  C_38_S_1_L_3_out, I4 =>  C_38_S_1_L_4_out, I5 =>  C_38_S_1_L_5_out); 
C_38_S_2_inst : LUT6 generic map(INIT => "1111111011101010111111101110100011101000100000001010100010000000") port map( O =>C_38_S_2_out, I0 =>  C_38_S_2_L_0_out, I1 =>  C_38_S_2_L_1_out, I2 =>  C_38_S_2_L_2_out, I3 =>  C_38_S_2_L_3_out, I4 =>  C_38_S_2_L_4_out, I5 =>  C_38_S_2_L_5_out); 
C_38_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001000100011101110111010001110100010000000") port map( O =>C_38_S_3_out, I0 =>  C_38_S_3_L_0_out, I1 =>  C_38_S_3_L_1_out, I2 =>  C_38_S_3_L_2_out, I3 =>  C_38_S_3_L_3_out, I4 =>  C_38_S_3_L_4_out, I5 =>  C_38_S_3_L_5_out); 
C_38_S_4_inst : LUT6 generic map(INIT => "1111111011101000111110101010000011111010101000001110100010000000") port map( O =>C_38_S_4_out, I0 =>  C_38_S_4_L_0_out, I1 =>  C_38_S_4_L_1_out, I2 =>  C_38_S_4_L_2_out, I3 =>  C_38_S_4_L_3_out, I4 =>  C_38_S_4_L_4_out, I5 =>  C_38_S_4_L_5_out); 
C_38_S_5_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_38_S_5_out, I0 =>  C_38_S_5_L_0_out, I1 =>  C_38_S_5_L_1_out, I2 =>  C_38_S_5_L_2_out, I3 =>  C_38_S_5_L_3_out, I4 =>  C_38_S_5_L_4_out, I5 =>  C_38_S_5_L_5_out); 

C_38_inst : LUT6 generic map(INIT => "1110101010101010101010101010100011101010101010101010101010101000") port map( O =>C_38_out, I0 =>  C_38_S_0_out, I1 =>  C_38_S_1_out, I2 =>  C_38_S_2_out, I3 =>  C_38_S_3_out, I4 =>  C_38_S_4_out, I5 =>  C_38_S_5_out); 

 
C_39_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_39_S_0_out, I0 =>  C_39_S_0_L_0_out, I1 =>  C_39_S_0_L_1_out, I2 =>  C_39_S_0_L_2_out, I3 =>  C_39_S_0_L_3_out, I4 =>  C_39_S_0_L_4_out, I5 =>  C_39_S_0_L_5_out); 
C_39_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_39_S_1_out, I0 =>  C_39_S_1_L_0_out, I1 =>  C_39_S_1_L_1_out, I2 =>  C_39_S_1_L_2_out, I3 =>  C_39_S_1_L_3_out, I4 =>  C_39_S_1_L_4_out, I5 =>  C_39_S_1_L_5_out); 
C_39_S_2_inst : LUT6 generic map(INIT => "1111111011101000111111001110100011101000110000001110100010000000") port map( O =>C_39_S_2_out, I0 =>  C_39_S_2_L_0_out, I1 =>  C_39_S_2_L_1_out, I2 =>  C_39_S_2_L_2_out, I3 =>  C_39_S_2_L_3_out, I4 =>  C_39_S_2_L_4_out, I5 =>  C_39_S_2_L_5_out); 
C_39_S_3_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_39_S_3_out, I0 =>  C_39_S_3_L_0_out, I1 =>  C_39_S_3_L_1_out, I2 =>  C_39_S_3_L_2_out, I3 =>  C_39_S_3_L_3_out, I4 =>  C_39_S_3_L_4_out, I5 =>  C_39_S_3_L_5_out); 
C_39_S_4_inst : LUT6 generic map(INIT => "1111111111111110111011101110100011101000100010001000000000000000") port map( O =>C_39_S_4_out, I0 =>  C_39_S_4_L_0_out, I1 =>  C_39_S_4_L_1_out, I2 =>  C_39_S_4_L_2_out, I3 =>  C_39_S_4_L_3_out, I4 =>  C_39_S_4_L_4_out, I5 =>  C_39_S_4_L_5_out); 
C_39_S_5_inst : LUT6 generic map(INIT => "1111111011101100111011001000100011101110110010001100100010000000") port map( O =>C_39_S_5_out, I0 =>  C_39_S_5_L_0_out, I1 =>  C_39_S_5_L_1_out, I2 =>  C_39_S_5_L_2_out, I3 =>  C_39_S_5_L_3_out, I4 =>  C_39_S_5_L_4_out, I5 =>  C_39_S_5_L_5_out); 

C_39_inst : LUT6 generic map(INIT => "1110101010101010111010101010101010101010101010001010101010101000") port map( O =>C_39_out, I0 =>  C_39_S_0_out, I1 =>  C_39_S_1_out, I2 =>  C_39_S_2_out, I3 =>  C_39_S_3_out, I4 =>  C_39_S_4_out, I5 =>  C_39_S_5_out); 

 
C_40_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_40_S_0_out, I0 =>  C_40_S_0_L_0_out, I1 =>  C_40_S_0_L_1_out, I2 =>  C_40_S_0_L_2_out, I3 =>  C_40_S_0_L_3_out, I4 =>  C_40_S_0_L_4_out, I5 =>  C_40_S_0_L_5_out); 
C_40_S_1_inst : LUT6 generic map(INIT => "1111111011101000111110101000000011111110101000001110100010000000") port map( O =>C_40_S_1_out, I0 =>  C_40_S_1_L_0_out, I1 =>  C_40_S_1_L_1_out, I2 =>  C_40_S_1_L_2_out, I3 =>  C_40_S_1_L_3_out, I4 =>  C_40_S_1_L_4_out, I5 =>  C_40_S_1_L_5_out); 
C_40_S_2_inst : LUT6 generic map(INIT => "1111111111101100111011101000100011101110100010001100100000000000") port map( O =>C_40_S_2_out, I0 =>  C_40_S_2_L_0_out, I1 =>  C_40_S_2_L_1_out, I2 =>  C_40_S_2_L_2_out, I3 =>  C_40_S_2_L_3_out, I4 =>  C_40_S_2_L_4_out, I5 =>  C_40_S_2_L_5_out); 
C_40_S_3_inst : LUT6 generic map(INIT => "1111111011101010111110101010100011101010101000001010100010000000") port map( O =>C_40_S_3_out, I0 =>  C_40_S_3_L_0_out, I1 =>  C_40_S_3_L_1_out, I2 =>  C_40_S_3_L_2_out, I3 =>  C_40_S_3_L_3_out, I4 =>  C_40_S_3_L_4_out, I5 =>  C_40_S_3_L_5_out); 
C_40_S_4_inst : LUT6 generic map(INIT => "1111111011101000111110101010000011111010101000001110100010000000") port map( O =>C_40_S_4_out, I0 =>  C_40_S_4_L_0_out, I1 =>  C_40_S_4_L_1_out, I2 =>  C_40_S_4_L_2_out, I3 =>  C_40_S_4_L_3_out, I4 =>  C_40_S_4_L_4_out, I5 =>  C_40_S_4_L_5_out); 
C_40_S_5_inst : LUT6 generic map(INIT => "1111111111101000111111101110100011101000100000001110100000000000") port map( O =>C_40_S_5_out, I0 =>  C_40_S_5_L_0_out, I1 =>  C_40_S_5_L_1_out, I2 =>  C_40_S_5_L_2_out, I3 =>  C_40_S_5_L_3_out, I4 =>  C_40_S_5_L_4_out, I5 =>  C_40_S_5_L_5_out); 

C_40_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_40_out, I0 =>  C_40_S_0_out, I1 =>  C_40_S_1_out, I2 =>  C_40_S_2_out, I3 =>  C_40_S_3_out, I4 =>  C_40_S_4_out, I5 =>  C_40_S_5_out); 

 
C_41_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_41_S_0_out, I0 =>  C_41_S_0_L_0_out, I1 =>  C_41_S_0_L_1_out, I2 =>  C_41_S_0_L_2_out, I3 =>  C_41_S_0_L_3_out, I4 =>  C_41_S_0_L_4_out, I5 =>  C_41_S_0_L_5_out); 
C_41_S_1_inst : LUT6 generic map(INIT => "1111111011101100111011101000100011101110100010001100100010000000") port map( O =>C_41_S_1_out, I0 =>  C_41_S_1_L_0_out, I1 =>  C_41_S_1_L_1_out, I2 =>  C_41_S_1_L_2_out, I3 =>  C_41_S_1_L_3_out, I4 =>  C_41_S_1_L_4_out, I5 =>  C_41_S_1_L_5_out); 
C_41_S_2_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_41_S_2_out, I0 =>  C_41_S_2_L_0_out, I1 =>  C_41_S_2_L_1_out, I2 =>  C_41_S_2_L_2_out, I3 =>  C_41_S_2_L_3_out, I4 =>  C_41_S_2_L_4_out, I5 =>  C_41_S_2_L_5_out); 
C_41_S_3_inst : LUT6 generic map(INIT => "1111111011111110111010001110100011101000111010001000000010000000") port map( O =>C_41_S_3_out, I0 =>  C_41_S_3_L_0_out, I1 =>  C_41_S_3_L_1_out, I2 =>  C_41_S_3_L_2_out, I3 =>  C_41_S_3_L_3_out, I4 =>  C_41_S_3_L_4_out, I5 =>  C_41_S_3_L_5_out); 
C_41_S_4_inst : LUT6 generic map(INIT => "1111111111101010111011101000000011111110100010001010100000000000") port map( O =>C_41_S_4_out, I0 =>  C_41_S_4_L_0_out, I1 =>  C_41_S_4_L_1_out, I2 =>  C_41_S_4_L_2_out, I3 =>  C_41_S_4_L_3_out, I4 =>  C_41_S_4_L_4_out, I5 =>  C_41_S_4_L_5_out); 
C_41_S_5_inst : LUT6 generic map(INIT => "1111111111111000111111101110000011111000100000001110000000000000") port map( O =>C_41_S_5_out, I0 =>  C_41_S_5_L_0_out, I1 =>  C_41_S_5_L_1_out, I2 =>  C_41_S_5_L_2_out, I3 =>  C_41_S_5_L_3_out, I4 =>  C_41_S_5_L_4_out, I5 =>  C_41_S_5_L_5_out); 

C_41_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_41_out, I0 =>  C_41_S_0_out, I1 =>  C_41_S_1_out, I2 =>  C_41_S_2_out, I3 =>  C_41_S_3_out, I4 =>  C_41_S_4_out, I5 =>  C_41_S_5_out); 

 
C_42_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010100011101010101010101010101010101000") port map( O =>C_42_S_0_out, I0 =>  C_42_S_0_L_0_out, I1 =>  C_42_S_0_L_1_out, I2 =>  C_42_S_0_L_2_out, I3 =>  C_42_S_0_L_3_out, I4 =>  C_42_S_0_L_4_out, I5 =>  C_42_S_0_L_5_out); 
C_42_S_1_inst : LUT6 generic map(INIT => "1110111011101000111011101110100011101000100010001110100010001000") port map( O =>C_42_S_1_out, I0 =>  C_42_S_1_L_0_out, I1 =>  C_42_S_1_L_1_out, I2 =>  C_42_S_1_L_2_out, I3 =>  C_42_S_1_L_3_out, I4 =>  C_42_S_1_L_4_out, I5 =>  C_42_S_1_L_5_out); 
C_42_S_2_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_42_S_2_out, I0 =>  C_42_S_2_L_0_out, I1 =>  C_42_S_2_L_1_out, I2 =>  C_42_S_2_L_2_out, I3 =>  C_42_S_2_L_3_out, I4 =>  C_42_S_2_L_4_out, I5 =>  C_42_S_2_L_5_out); 
C_42_S_3_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_42_S_3_out, I0 =>  C_42_S_3_L_0_out, I1 =>  C_42_S_3_L_1_out, I2 =>  C_42_S_3_L_2_out, I3 =>  C_42_S_3_L_3_out, I4 =>  C_42_S_3_L_4_out, I5 =>  C_42_S_3_L_5_out); 
C_42_S_4_inst : LUT6 generic map(INIT => "1111111011101000111010101110100011101000101010001110100010000000") port map( O =>C_42_S_4_out, I0 =>  C_42_S_4_L_0_out, I1 =>  C_42_S_4_L_1_out, I2 =>  C_42_S_4_L_2_out, I3 =>  C_42_S_4_L_3_out, I4 =>  C_42_S_4_L_4_out, I5 =>  C_42_S_4_L_5_out); 
C_42_S_5_inst : LUT6 generic map(INIT => "1111111011111110111010001010000011111010111010001000000010000000") port map( O =>C_42_S_5_out, I0 =>  C_42_S_5_L_0_out, I1 =>  C_42_S_5_L_1_out, I2 =>  C_42_S_5_L_2_out, I3 =>  C_42_S_5_L_3_out, I4 =>  C_42_S_5_L_4_out, I5 =>  C_42_S_5_L_5_out); 

C_42_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_42_out, I0 =>  C_42_S_0_out, I1 =>  C_42_S_1_out, I2 =>  C_42_S_2_out, I3 =>  C_42_S_3_out, I4 =>  C_42_S_4_out, I5 =>  C_42_S_5_out); 

 
C_43_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_43_S_0_out, I0 =>  C_43_S_0_L_0_out, I1 =>  C_43_S_0_L_1_out, I2 =>  C_43_S_0_L_2_out, I3 =>  C_43_S_0_L_3_out, I4 =>  C_43_S_0_L_4_out, I5 =>  C_43_S_0_L_5_out); 
C_43_S_1_inst : LUT6 generic map(INIT => "1110101010101010111010101010100011101010101010001010101010101000") port map( O =>C_43_S_1_out, I0 =>  C_43_S_1_L_0_out, I1 =>  C_43_S_1_L_1_out, I2 =>  C_43_S_1_L_2_out, I3 =>  C_43_S_1_L_3_out, I4 =>  C_43_S_1_L_4_out, I5 =>  C_43_S_1_L_5_out); 
C_43_S_2_inst : LUT6 generic map(INIT => "1111111011101000111111001100000011111100110000001110100010000000") port map( O =>C_43_S_2_out, I0 =>  C_43_S_2_L_0_out, I1 =>  C_43_S_2_L_1_out, I2 =>  C_43_S_2_L_2_out, I3 =>  C_43_S_2_L_3_out, I4 =>  C_43_S_2_L_4_out, I5 =>  C_43_S_2_L_5_out); 
C_43_S_3_inst : LUT6 generic map(INIT => "1111111111111110111010101010100011101010101010001000000000000000") port map( O =>C_43_S_3_out, I0 =>  C_43_S_3_L_0_out, I1 =>  C_43_S_3_L_1_out, I2 =>  C_43_S_3_L_2_out, I3 =>  C_43_S_3_L_3_out, I4 =>  C_43_S_3_L_4_out, I5 =>  C_43_S_3_L_5_out); 
C_43_S_4_inst : LUT6 generic map(INIT => "1111111011101000111110001110000011111000111000001110100010000000") port map( O =>C_43_S_4_out, I0 =>  C_43_S_4_L_0_out, I1 =>  C_43_S_4_L_1_out, I2 =>  C_43_S_4_L_2_out, I3 =>  C_43_S_4_L_3_out, I4 =>  C_43_S_4_L_4_out, I5 =>  C_43_S_4_L_5_out); 
C_43_S_5_inst : LUT6 generic map(INIT => "1111111011111100111111001110100011101000110000001100000010000000") port map( O =>C_43_S_5_out, I0 =>  C_43_S_5_L_0_out, I1 =>  C_43_S_5_L_1_out, I2 =>  C_43_S_5_L_2_out, I3 =>  C_43_S_5_L_3_out, I4 =>  C_43_S_5_L_4_out, I5 =>  C_43_S_5_L_5_out); 

C_43_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_43_out, I0 =>  C_43_S_0_out, I1 =>  C_43_S_1_out, I2 =>  C_43_S_2_out, I3 =>  C_43_S_3_out, I4 =>  C_43_S_4_out, I5 =>  C_43_S_5_out); 

 
C_44_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_44_S_0_out, I0 =>  C_44_S_0_L_0_out, I1 =>  C_44_S_0_L_1_out, I2 =>  C_44_S_0_L_2_out, I3 =>  C_44_S_0_L_3_out, I4 =>  C_44_S_0_L_4_out, I5 =>  C_44_S_0_L_5_out); 
C_44_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_44_S_1_out, I0 =>  C_44_S_1_L_0_out, I1 =>  C_44_S_1_L_1_out, I2 =>  C_44_S_1_L_2_out, I3 =>  C_44_S_1_L_3_out, I4 =>  C_44_S_1_L_4_out, I5 =>  C_44_S_1_L_5_out); 
C_44_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010101010000011111010101010001110100010000000") port map( O =>C_44_S_2_out, I0 =>  C_44_S_2_L_0_out, I1 =>  C_44_S_2_L_1_out, I2 =>  C_44_S_2_L_2_out, I3 =>  C_44_S_2_L_3_out, I4 =>  C_44_S_2_L_4_out, I5 =>  C_44_S_2_L_5_out); 
C_44_S_3_inst : LUT6 generic map(INIT => "1111111111111110111010001000000011111110111010001000000000000000") port map( O =>C_44_S_3_out, I0 =>  C_44_S_3_L_0_out, I1 =>  C_44_S_3_L_1_out, I2 =>  C_44_S_3_L_2_out, I3 =>  C_44_S_3_L_3_out, I4 =>  C_44_S_3_L_4_out, I5 =>  C_44_S_3_L_5_out); 
C_44_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_44_S_4_out, I0 =>  C_44_S_4_L_0_out, I1 =>  C_44_S_4_L_1_out, I2 =>  C_44_S_4_L_2_out, I3 =>  C_44_S_4_L_3_out, I4 =>  C_44_S_4_L_4_out, I5 =>  C_44_S_4_L_5_out); 
C_44_S_5_inst : LUT6 generic map(INIT => "1111111011101010111110101110100011101000101000001010100010000000") port map( O =>C_44_S_5_out, I0 =>  C_44_S_5_L_0_out, I1 =>  C_44_S_5_L_1_out, I2 =>  C_44_S_5_L_2_out, I3 =>  C_44_S_5_L_3_out, I4 =>  C_44_S_5_L_4_out, I5 =>  C_44_S_5_L_5_out); 

C_44_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_44_out, I0 =>  C_44_S_0_out, I1 =>  C_44_S_1_out, I2 =>  C_44_S_2_out, I3 =>  C_44_S_3_out, I4 =>  C_44_S_4_out, I5 =>  C_44_S_5_out); 

 
C_45_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_45_S_0_out, I0 =>  C_45_S_0_L_0_out, I1 =>  C_45_S_0_L_1_out, I2 =>  C_45_S_0_L_2_out, I3 =>  C_45_S_0_L_3_out, I4 =>  C_45_S_0_L_4_out, I5 =>  C_45_S_0_L_5_out); 
C_45_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010001010100011101010111010001010100010000000") port map( O =>C_45_S_1_out, I0 =>  C_45_S_1_L_0_out, I1 =>  C_45_S_1_L_1_out, I2 =>  C_45_S_1_L_2_out, I3 =>  C_45_S_1_L_3_out, I4 =>  C_45_S_1_L_4_out, I5 =>  C_45_S_1_L_5_out); 
C_45_S_2_inst : LUT6 generic map(INIT => "1111111011101010111011101010100011101010100010001010100010000000") port map( O =>C_45_S_2_out, I0 =>  C_45_S_2_L_0_out, I1 =>  C_45_S_2_L_1_out, I2 =>  C_45_S_2_L_2_out, I3 =>  C_45_S_2_L_3_out, I4 =>  C_45_S_2_L_4_out, I5 =>  C_45_S_2_L_5_out); 
C_45_S_3_inst : LUT6 generic map(INIT => "1111111111101000111111101110000011111000100000001110100000000000") port map( O =>C_45_S_3_out, I0 =>  C_45_S_3_L_0_out, I1 =>  C_45_S_3_L_1_out, I2 =>  C_45_S_3_L_2_out, I3 =>  C_45_S_3_L_3_out, I4 =>  C_45_S_3_L_4_out, I5 =>  C_45_S_3_L_5_out); 
C_45_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_45_S_4_out, I0 =>  C_45_S_4_L_0_out, I1 =>  C_45_S_4_L_1_out, I2 =>  C_45_S_4_L_2_out, I3 =>  C_45_S_4_L_3_out, I4 =>  C_45_S_4_L_4_out, I5 =>  C_45_S_4_L_5_out); 
C_45_S_5_inst : LUT6 generic map(INIT => "1111111111101000111111101000000011111110100000001110100000000000") port map( O =>C_45_S_5_out, I0 =>  C_45_S_5_L_0_out, I1 =>  C_45_S_5_L_1_out, I2 =>  C_45_S_5_L_2_out, I3 =>  C_45_S_5_L_3_out, I4 =>  C_45_S_5_L_4_out, I5 =>  C_45_S_5_L_5_out); 

C_45_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_45_out, I0 =>  C_45_S_0_out, I1 =>  C_45_S_1_out, I2 =>  C_45_S_2_out, I3 =>  C_45_S_3_out, I4 =>  C_45_S_4_out, I5 =>  C_45_S_5_out); 

 
C_46_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_46_S_0_out, I0 =>  C_46_S_0_L_0_out, I1 =>  C_46_S_0_L_1_out, I2 =>  C_46_S_0_L_2_out, I3 =>  C_46_S_0_L_3_out, I4 =>  C_46_S_0_L_4_out, I5 =>  C_46_S_0_L_5_out); 
C_46_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_46_S_1_out, I0 =>  C_46_S_1_L_0_out, I1 =>  C_46_S_1_L_1_out, I2 =>  C_46_S_1_L_2_out, I3 =>  C_46_S_1_L_3_out, I4 =>  C_46_S_1_L_4_out, I5 =>  C_46_S_1_L_5_out); 
C_46_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101110100011101000101010001010100010000000") port map( O =>C_46_S_2_out, I0 =>  C_46_S_2_L_0_out, I1 =>  C_46_S_2_L_1_out, I2 =>  C_46_S_2_L_2_out, I3 =>  C_46_S_2_L_3_out, I4 =>  C_46_S_2_L_4_out, I5 =>  C_46_S_2_L_5_out); 
C_46_S_3_inst : LUT6 generic map(INIT => "1111111111111110111011101100100011101100100010001000000000000000") port map( O =>C_46_S_3_out, I0 =>  C_46_S_3_L_0_out, I1 =>  C_46_S_3_L_1_out, I2 =>  C_46_S_3_L_2_out, I3 =>  C_46_S_3_L_3_out, I4 =>  C_46_S_3_L_4_out, I5 =>  C_46_S_3_L_5_out); 
C_46_S_4_inst : LUT6 generic map(INIT => "1111111011101000111010001110000011111000111010001110100010000000") port map( O =>C_46_S_4_out, I0 =>  C_46_S_4_L_0_out, I1 =>  C_46_S_4_L_1_out, I2 =>  C_46_S_4_L_2_out, I3 =>  C_46_S_4_L_3_out, I4 =>  C_46_S_4_L_4_out, I5 =>  C_46_S_4_L_5_out); 
C_46_S_5_inst : LUT6 generic map(INIT => "1111111011111000111110001110100011101000111000001110000010000000") port map( O =>C_46_S_5_out, I0 =>  C_46_S_5_L_0_out, I1 =>  C_46_S_5_L_1_out, I2 =>  C_46_S_5_L_2_out, I3 =>  C_46_S_5_L_3_out, I4 =>  C_46_S_5_L_4_out, I5 =>  C_46_S_5_L_5_out); 

C_46_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_46_out, I0 =>  C_46_S_0_out, I1 =>  C_46_S_1_out, I2 =>  C_46_S_2_out, I3 =>  C_46_S_3_out, I4 =>  C_46_S_4_out, I5 =>  C_46_S_5_out); 

 
C_47_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_47_S_0_out, I0 =>  C_47_S_0_L_0_out, I1 =>  C_47_S_0_L_1_out, I2 =>  C_47_S_0_L_2_out, I3 =>  C_47_S_0_L_3_out, I4 =>  C_47_S_0_L_4_out, I5 =>  C_47_S_0_L_5_out); 
C_47_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010001000100011101110111010001110100010000000") port map( O =>C_47_S_1_out, I0 =>  C_47_S_1_L_0_out, I1 =>  C_47_S_1_L_1_out, I2 =>  C_47_S_1_L_2_out, I3 =>  C_47_S_1_L_3_out, I4 =>  C_47_S_1_L_4_out, I5 =>  C_47_S_1_L_5_out); 
C_47_S_2_inst : LUT6 generic map(INIT => "1111111111111110111010001000000011111110111010001000000000000000") port map( O =>C_47_S_2_out, I0 =>  C_47_S_2_L_0_out, I1 =>  C_47_S_2_L_1_out, I2 =>  C_47_S_2_L_2_out, I3 =>  C_47_S_2_L_3_out, I4 =>  C_47_S_2_L_4_out, I5 =>  C_47_S_2_L_5_out); 
C_47_S_3_inst : LUT6 generic map(INIT => "1111111111111000111111001110000011111000110000001110000000000000") port map( O =>C_47_S_3_out, I0 =>  C_47_S_3_L_0_out, I1 =>  C_47_S_3_L_1_out, I2 =>  C_47_S_3_L_2_out, I3 =>  C_47_S_3_L_3_out, I4 =>  C_47_S_3_L_4_out, I5 =>  C_47_S_3_L_5_out); 
C_47_S_4_inst : LUT6 generic map(INIT => "1111111011101100111111101110100011101000100000001100100010000000") port map( O =>C_47_S_4_out, I0 =>  C_47_S_4_L_0_out, I1 =>  C_47_S_4_L_1_out, I2 =>  C_47_S_4_L_2_out, I3 =>  C_47_S_4_L_3_out, I4 =>  C_47_S_4_L_4_out, I5 =>  C_47_S_4_L_5_out); 
C_47_S_5_inst : LUT6 generic map(INIT => "1111111111101000111111101010100011101010100000001110100000000000") port map( O =>C_47_S_5_out, I0 =>  C_47_S_5_L_0_out, I1 =>  C_47_S_5_L_1_out, I2 =>  C_47_S_5_L_2_out, I3 =>  C_47_S_5_L_3_out, I4 =>  C_47_S_5_L_4_out, I5 =>  C_47_S_5_L_5_out); 

C_47_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_47_out, I0 =>  C_47_S_0_out, I1 =>  C_47_S_1_out, I2 =>  C_47_S_2_out, I3 =>  C_47_S_3_out, I4 =>  C_47_S_4_out, I5 =>  C_47_S_5_out); 

 
C_48_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_48_S_0_out, I0 =>  C_48_S_0_L_0_out, I1 =>  C_48_S_0_L_1_out, I2 =>  C_48_S_0_L_2_out, I3 =>  C_48_S_0_L_3_out, I4 =>  C_48_S_0_L_4_out, I5 =>  C_48_S_0_L_5_out); 
C_48_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_48_S_1_out, I0 =>  C_48_S_1_L_0_out, I1 =>  C_48_S_1_L_1_out, I2 =>  C_48_S_1_L_2_out, I3 =>  C_48_S_1_L_3_out, I4 =>  C_48_S_1_L_4_out, I5 =>  C_48_S_1_L_5_out); 
C_48_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_48_S_2_out, I0 =>  C_48_S_2_L_0_out, I1 =>  C_48_S_2_L_1_out, I2 =>  C_48_S_2_L_2_out, I3 =>  C_48_S_2_L_3_out, I4 =>  C_48_S_2_L_4_out, I5 =>  C_48_S_2_L_5_out); 
C_48_S_3_inst : LUT6 generic map(INIT => "1111111111111010111110001110000011111000111000001010000000000000") port map( O =>C_48_S_3_out, I0 =>  C_48_S_3_L_0_out, I1 =>  C_48_S_3_L_1_out, I2 =>  C_48_S_3_L_2_out, I3 =>  C_48_S_3_L_3_out, I4 =>  C_48_S_3_L_4_out, I5 =>  C_48_S_3_L_5_out); 
C_48_S_4_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_48_S_4_out, I0 =>  C_48_S_4_L_0_out, I1 =>  C_48_S_4_L_1_out, I2 =>  C_48_S_4_L_2_out, I3 =>  C_48_S_4_L_3_out, I4 =>  C_48_S_4_L_4_out, I5 =>  C_48_S_4_L_5_out); 
C_48_S_5_inst : LUT6 generic map(INIT => "1111111111101010111010101010000011111010101010001010100000000000") port map( O =>C_48_S_5_out, I0 =>  C_48_S_5_L_0_out, I1 =>  C_48_S_5_L_1_out, I2 =>  C_48_S_5_L_2_out, I3 =>  C_48_S_5_L_3_out, I4 =>  C_48_S_5_L_4_out, I5 =>  C_48_S_5_L_5_out); 

C_48_inst : LUT6 generic map(INIT => "1110101010101010111010101010100011101010101010001010101010101000") port map( O =>C_48_out, I0 =>  C_48_S_0_out, I1 =>  C_48_S_1_out, I2 =>  C_48_S_2_out, I3 =>  C_48_S_3_out, I4 =>  C_48_S_4_out, I5 =>  C_48_S_5_out); 

 
C_49_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_49_S_0_out, I0 =>  C_49_S_0_L_0_out, I1 =>  C_49_S_0_L_1_out, I2 =>  C_49_S_0_L_2_out, I3 =>  C_49_S_0_L_3_out, I4 =>  C_49_S_0_L_4_out, I5 =>  C_49_S_0_L_5_out); 
C_49_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010001010100011101010111010001010100010000000") port map( O =>C_49_S_1_out, I0 =>  C_49_S_1_L_0_out, I1 =>  C_49_S_1_L_1_out, I2 =>  C_49_S_1_L_2_out, I3 =>  C_49_S_1_L_3_out, I4 =>  C_49_S_1_L_4_out, I5 =>  C_49_S_1_L_5_out); 
C_49_S_2_inst : LUT6 generic map(INIT => "1111111011101100111011001110100011101000110010001100100010000000") port map( O =>C_49_S_2_out, I0 =>  C_49_S_2_L_0_out, I1 =>  C_49_S_2_L_1_out, I2 =>  C_49_S_2_L_2_out, I3 =>  C_49_S_2_L_3_out, I4 =>  C_49_S_2_L_4_out, I5 =>  C_49_S_2_L_5_out); 
C_49_S_3_inst : LUT6 generic map(INIT => "1111111011111110111011101110100011101000100010001000000010000000") port map( O =>C_49_S_3_out, I0 =>  C_49_S_3_L_0_out, I1 =>  C_49_S_3_L_1_out, I2 =>  C_49_S_3_L_2_out, I3 =>  C_49_S_3_L_3_out, I4 =>  C_49_S_3_L_4_out, I5 =>  C_49_S_3_L_5_out); 
C_49_S_4_inst : LUT6 generic map(INIT => "1111111011101000111011101000100011101110100010001110100010000000") port map( O =>C_49_S_4_out, I0 =>  C_49_S_4_L_0_out, I1 =>  C_49_S_4_L_1_out, I2 =>  C_49_S_4_L_2_out, I3 =>  C_49_S_4_L_3_out, I4 =>  C_49_S_4_L_4_out, I5 =>  C_49_S_4_L_5_out); 
C_49_S_5_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_49_S_5_out, I0 =>  C_49_S_5_L_0_out, I1 =>  C_49_S_5_L_1_out, I2 =>  C_49_S_5_L_2_out, I3 =>  C_49_S_5_L_3_out, I4 =>  C_49_S_5_L_4_out, I5 =>  C_49_S_5_L_5_out); 

C_49_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_49_out, I0 =>  C_49_S_0_out, I1 =>  C_49_S_1_out, I2 =>  C_49_S_2_out, I3 =>  C_49_S_3_out, I4 =>  C_49_S_4_out, I5 =>  C_49_S_5_out); 

 
C_50_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_50_S_0_out, I0 =>  C_50_S_0_L_0_out, I1 =>  C_50_S_0_L_1_out, I2 =>  C_50_S_0_L_2_out, I3 =>  C_50_S_0_L_3_out, I4 =>  C_50_S_0_L_4_out, I5 =>  C_50_S_0_L_5_out); 
C_50_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_50_S_1_out, I0 =>  C_50_S_1_L_0_out, I1 =>  C_50_S_1_L_1_out, I2 =>  C_50_S_1_L_2_out, I3 =>  C_50_S_1_L_3_out, I4 =>  C_50_S_1_L_4_out, I5 =>  C_50_S_1_L_5_out); 
C_50_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001110000011111000111010001110100010000000") port map( O =>C_50_S_2_out, I0 =>  C_50_S_2_L_0_out, I1 =>  C_50_S_2_L_1_out, I2 =>  C_50_S_2_L_2_out, I3 =>  C_50_S_2_L_3_out, I4 =>  C_50_S_2_L_4_out, I5 =>  C_50_S_2_L_5_out); 
C_50_S_3_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_50_S_3_out, I0 =>  C_50_S_3_L_0_out, I1 =>  C_50_S_3_L_1_out, I2 =>  C_50_S_3_L_2_out, I3 =>  C_50_S_3_L_3_out, I4 =>  C_50_S_3_L_4_out, I5 =>  C_50_S_3_L_5_out); 
C_50_S_4_inst : LUT6 generic map(INIT => "1111111011111110111010001010100011101010111010001000000010000000") port map( O =>C_50_S_4_out, I0 =>  C_50_S_4_L_0_out, I1 =>  C_50_S_4_L_1_out, I2 =>  C_50_S_4_L_2_out, I3 =>  C_50_S_4_L_3_out, I4 =>  C_50_S_4_L_4_out, I5 =>  C_50_S_4_L_5_out); 
C_50_S_5_inst : LUT6 generic map(INIT => "1111111011101100111010001000000011111110111010001100100010000000") port map( O =>C_50_S_5_out, I0 =>  C_50_S_5_L_0_out, I1 =>  C_50_S_5_L_1_out, I2 =>  C_50_S_5_L_2_out, I3 =>  C_50_S_5_L_3_out, I4 =>  C_50_S_5_L_4_out, I5 =>  C_50_S_5_L_5_out); 

C_50_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_50_out, I0 =>  C_50_S_0_out, I1 =>  C_50_S_1_out, I2 =>  C_50_S_2_out, I3 =>  C_50_S_3_out, I4 =>  C_50_S_4_out, I5 =>  C_50_S_5_out); 

 
C_51_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_51_S_0_out, I0 =>  C_51_S_0_L_0_out, I1 =>  C_51_S_0_L_1_out, I2 =>  C_51_S_0_L_2_out, I3 =>  C_51_S_0_L_3_out, I4 =>  C_51_S_0_L_4_out, I5 =>  C_51_S_0_L_5_out); 
C_51_S_1_inst : LUT6 generic map(INIT => "1111111011101110111010001110100011101000111010001000100010000000") port map( O =>C_51_S_1_out, I0 =>  C_51_S_1_L_0_out, I1 =>  C_51_S_1_L_1_out, I2 =>  C_51_S_1_L_2_out, I3 =>  C_51_S_1_L_3_out, I4 =>  C_51_S_1_L_4_out, I5 =>  C_51_S_1_L_5_out); 
C_51_S_2_inst : LUT6 generic map(INIT => "1111111011111000111110001100000011111100111000001110000010000000") port map( O =>C_51_S_2_out, I0 =>  C_51_S_2_L_0_out, I1 =>  C_51_S_2_L_1_out, I2 =>  C_51_S_2_L_2_out, I3 =>  C_51_S_2_L_3_out, I4 =>  C_51_S_2_L_4_out, I5 =>  C_51_S_2_L_5_out); 
C_51_S_3_inst : LUT6 generic map(INIT => "1111111011101100111010001000100011101110111010001100100010000000") port map( O =>C_51_S_3_out, I0 =>  C_51_S_3_L_0_out, I1 =>  C_51_S_3_L_1_out, I2 =>  C_51_S_3_L_2_out, I3 =>  C_51_S_3_L_3_out, I4 =>  C_51_S_3_L_4_out, I5 =>  C_51_S_3_L_5_out); 
C_51_S_4_inst : LUT6 generic map(INIT => "1111111011111110111010001110100011101000111010001000000010000000") port map( O =>C_51_S_4_out, I0 =>  C_51_S_4_L_0_out, I1 =>  C_51_S_4_L_1_out, I2 =>  C_51_S_4_L_2_out, I3 =>  C_51_S_4_L_3_out, I4 =>  C_51_S_4_L_4_out, I5 =>  C_51_S_4_L_5_out); 
C_51_S_5_inst : LUT6 generic map(INIT => "1111111111111110111010001000000011111110111010001000000000000000") port map( O =>C_51_S_5_out, I0 =>  C_51_S_5_L_0_out, I1 =>  C_51_S_5_L_1_out, I2 =>  C_51_S_5_L_2_out, I3 =>  C_51_S_5_L_3_out, I4 =>  C_51_S_5_L_4_out, I5 =>  C_51_S_5_L_5_out); 

C_51_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_51_out, I0 =>  C_51_S_0_out, I1 =>  C_51_S_1_out, I2 =>  C_51_S_2_out, I3 =>  C_51_S_3_out, I4 =>  C_51_S_4_out, I5 =>  C_51_S_5_out); 

 
C_52_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_52_S_0_out, I0 =>  C_52_S_0_L_0_out, I1 =>  C_52_S_0_L_1_out, I2 =>  C_52_S_0_L_2_out, I3 =>  C_52_S_0_L_3_out, I4 =>  C_52_S_0_L_4_out, I5 =>  C_52_S_0_L_5_out); 
C_52_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_52_S_1_out, I0 =>  C_52_S_1_L_0_out, I1 =>  C_52_S_1_L_1_out, I2 =>  C_52_S_1_L_2_out, I3 =>  C_52_S_1_L_3_out, I4 =>  C_52_S_1_L_4_out, I5 =>  C_52_S_1_L_5_out); 
C_52_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_52_S_2_out, I0 =>  C_52_S_2_L_0_out, I1 =>  C_52_S_2_L_1_out, I2 =>  C_52_S_2_L_2_out, I3 =>  C_52_S_2_L_3_out, I4 =>  C_52_S_2_L_4_out, I5 =>  C_52_S_2_L_5_out); 
C_52_S_3_inst : LUT6 generic map(INIT => "1111111111111110111110101010100011101010101000001000000000000000") port map( O =>C_52_S_3_out, I0 =>  C_52_S_3_L_0_out, I1 =>  C_52_S_3_L_1_out, I2 =>  C_52_S_3_L_2_out, I3 =>  C_52_S_3_L_3_out, I4 =>  C_52_S_3_L_4_out, I5 =>  C_52_S_3_L_5_out); 
C_52_S_4_inst : LUT6 generic map(INIT => "1111111111101110111011101000100011101110100010001000100000000000") port map( O =>C_52_S_4_out, I0 =>  C_52_S_4_L_0_out, I1 =>  C_52_S_4_L_1_out, I2 =>  C_52_S_4_L_2_out, I3 =>  C_52_S_4_L_3_out, I4 =>  C_52_S_4_L_4_out, I5 =>  C_52_S_4_L_5_out); 
C_52_S_5_inst : LUT6 generic map(INIT => "1111111111101010111111101000100011101110100000001010100000000000") port map( O =>C_52_S_5_out, I0 =>  C_52_S_5_L_0_out, I1 =>  C_52_S_5_L_1_out, I2 =>  C_52_S_5_L_2_out, I3 =>  C_52_S_5_L_3_out, I4 =>  C_52_S_5_L_4_out, I5 =>  C_52_S_5_L_5_out); 

C_52_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_52_out, I0 =>  C_52_S_0_out, I1 =>  C_52_S_1_out, I2 =>  C_52_S_2_out, I3 =>  C_52_S_3_out, I4 =>  C_52_S_4_out, I5 =>  C_52_S_5_out); 

 
C_53_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_53_S_0_out, I0 =>  C_53_S_0_L_0_out, I1 =>  C_53_S_0_L_1_out, I2 =>  C_53_S_0_L_2_out, I3 =>  C_53_S_0_L_3_out, I4 =>  C_53_S_0_L_4_out, I5 =>  C_53_S_0_L_5_out); 
C_53_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_53_S_1_out, I0 =>  C_53_S_1_L_0_out, I1 =>  C_53_S_1_L_1_out, I2 =>  C_53_S_1_L_2_out, I3 =>  C_53_S_1_L_3_out, I4 =>  C_53_S_1_L_4_out, I5 =>  C_53_S_1_L_5_out); 
C_53_S_2_inst : LUT6 generic map(INIT => "1111111011101000111111101110100011101000100000001110100010000000") port map( O =>C_53_S_2_out, I0 =>  C_53_S_2_L_0_out, I1 =>  C_53_S_2_L_1_out, I2 =>  C_53_S_2_L_2_out, I3 =>  C_53_S_2_L_3_out, I4 =>  C_53_S_2_L_4_out, I5 =>  C_53_S_2_L_5_out); 
C_53_S_3_inst : LUT6 generic map(INIT => "1111111011101000111010001100100011101100111010001110100010000000") port map( O =>C_53_S_3_out, I0 =>  C_53_S_3_L_0_out, I1 =>  C_53_S_3_L_1_out, I2 =>  C_53_S_3_L_2_out, I3 =>  C_53_S_3_L_3_out, I4 =>  C_53_S_3_L_4_out, I5 =>  C_53_S_3_L_5_out); 
C_53_S_4_inst : LUT6 generic map(INIT => "1111111011111100111110001110000011111000111000001100000010000000") port map( O =>C_53_S_4_out, I0 =>  C_53_S_4_L_0_out, I1 =>  C_53_S_4_L_1_out, I2 =>  C_53_S_4_L_2_out, I3 =>  C_53_S_4_L_3_out, I4 =>  C_53_S_4_L_4_out, I5 =>  C_53_S_4_L_5_out); 
C_53_S_5_inst : LUT6 generic map(INIT => "1111111011101100111011001100100011101100110010001100100010000000") port map( O =>C_53_S_5_out, I0 =>  C_53_S_5_L_0_out, I1 =>  C_53_S_5_L_1_out, I2 =>  C_53_S_5_L_2_out, I3 =>  C_53_S_5_L_3_out, I4 =>  C_53_S_5_L_4_out, I5 =>  C_53_S_5_L_5_out); 

C_53_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_53_out, I0 =>  C_53_S_0_out, I1 =>  C_53_S_1_out, I2 =>  C_53_S_2_out, I3 =>  C_53_S_3_out, I4 =>  C_53_S_4_out, I5 =>  C_53_S_5_out); 

 
C_54_S_0_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_54_S_0_out, I0 =>  C_54_S_0_L_0_out, I1 =>  C_54_S_0_L_1_out, I2 =>  C_54_S_0_L_2_out, I3 =>  C_54_S_0_L_3_out, I4 =>  C_54_S_0_L_4_out, I5 =>  C_54_S_0_L_5_out); 
C_54_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_54_S_1_out, I0 =>  C_54_S_1_L_0_out, I1 =>  C_54_S_1_L_1_out, I2 =>  C_54_S_1_L_2_out, I3 =>  C_54_S_1_L_3_out, I4 =>  C_54_S_1_L_4_out, I5 =>  C_54_S_1_L_5_out); 
C_54_S_2_inst : LUT6 generic map(INIT => "1111111011101010111010001110100011101000111010001010100010000000") port map( O =>C_54_S_2_out, I0 =>  C_54_S_2_L_0_out, I1 =>  C_54_S_2_L_1_out, I2 =>  C_54_S_2_L_2_out, I3 =>  C_54_S_2_L_3_out, I4 =>  C_54_S_2_L_4_out, I5 =>  C_54_S_2_L_5_out); 
C_54_S_3_inst : LUT6 generic map(INIT => "1111111011101100111010001000000011111110111010001100100010000000") port map( O =>C_54_S_3_out, I0 =>  C_54_S_3_L_0_out, I1 =>  C_54_S_3_L_1_out, I2 =>  C_54_S_3_L_2_out, I3 =>  C_54_S_3_L_3_out, I4 =>  C_54_S_3_L_4_out, I5 =>  C_54_S_3_L_5_out); 
C_54_S_4_inst : LUT6 generic map(INIT => "1111111011101000111111101110000011111000100000001110100010000000") port map( O =>C_54_S_4_out, I0 =>  C_54_S_4_L_0_out, I1 =>  C_54_S_4_L_1_out, I2 =>  C_54_S_4_L_2_out, I3 =>  C_54_S_4_L_3_out, I4 =>  C_54_S_4_L_4_out, I5 =>  C_54_S_4_L_5_out); 
C_54_S_5_inst : LUT6 generic map(INIT => "1111111111111010111010101010100011101010101010001010000000000000") port map( O =>C_54_S_5_out, I0 =>  C_54_S_5_L_0_out, I1 =>  C_54_S_5_L_1_out, I2 =>  C_54_S_5_L_2_out, I3 =>  C_54_S_5_L_3_out, I4 =>  C_54_S_5_L_4_out, I5 =>  C_54_S_5_L_5_out); 

C_54_inst : LUT6 generic map(INIT => "1110101011101010111010101010100011101010101010001010100010101000") port map( O =>C_54_out, I0 =>  C_54_S_0_out, I1 =>  C_54_S_1_out, I2 =>  C_54_S_2_out, I3 =>  C_54_S_3_out, I4 =>  C_54_S_4_out, I5 =>  C_54_S_5_out); 

 
C_55_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_55_S_0_out, I0 =>  C_55_S_0_L_0_out, I1 =>  C_55_S_0_L_1_out, I2 =>  C_55_S_0_L_2_out, I3 =>  C_55_S_0_L_3_out, I4 =>  C_55_S_0_L_4_out, I5 =>  C_55_S_0_L_5_out); 
C_55_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_55_S_1_out, I0 =>  C_55_S_1_L_0_out, I1 =>  C_55_S_1_L_1_out, I2 =>  C_55_S_1_L_2_out, I3 =>  C_55_S_1_L_3_out, I4 =>  C_55_S_1_L_4_out, I5 =>  C_55_S_1_L_5_out); 
C_55_S_2_inst : LUT6 generic map(INIT => "1111111011111000111111101110000011111000100000001110000010000000") port map( O =>C_55_S_2_out, I0 =>  C_55_S_2_L_0_out, I1 =>  C_55_S_2_L_1_out, I2 =>  C_55_S_2_L_2_out, I3 =>  C_55_S_2_L_3_out, I4 =>  C_55_S_2_L_4_out, I5 =>  C_55_S_2_L_5_out); 
C_55_S_3_inst : LUT6 generic map(INIT => "1111111111101110111011101000100011101110100010001000100000000000") port map( O =>C_55_S_3_out, I0 =>  C_55_S_3_L_0_out, I1 =>  C_55_S_3_L_1_out, I2 =>  C_55_S_3_L_2_out, I3 =>  C_55_S_3_L_3_out, I4 =>  C_55_S_3_L_4_out, I5 =>  C_55_S_3_L_5_out); 
C_55_S_4_inst : LUT6 generic map(INIT => "1111111111101100111011001000100011101110110010001100100000000000") port map( O =>C_55_S_4_out, I0 =>  C_55_S_4_L_0_out, I1 =>  C_55_S_4_L_1_out, I2 =>  C_55_S_4_L_2_out, I3 =>  C_55_S_4_L_3_out, I4 =>  C_55_S_4_L_4_out, I5 =>  C_55_S_4_L_5_out); 
C_55_S_5_inst : LUT6 generic map(INIT => "1111111011111110111010001110000011111000111010001000000010000000") port map( O =>C_55_S_5_out, I0 =>  C_55_S_5_L_0_out, I1 =>  C_55_S_5_L_1_out, I2 =>  C_55_S_5_L_2_out, I3 =>  C_55_S_5_L_3_out, I4 =>  C_55_S_5_L_4_out, I5 =>  C_55_S_5_L_5_out); 

C_55_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_55_out, I0 =>  C_55_S_0_out, I1 =>  C_55_S_1_out, I2 =>  C_55_S_2_out, I3 =>  C_55_S_3_out, I4 =>  C_55_S_4_out, I5 =>  C_55_S_5_out); 

 
C_56_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_56_S_0_out, I0 =>  C_56_S_0_L_0_out, I1 =>  C_56_S_0_L_1_out, I2 =>  C_56_S_0_L_2_out, I3 =>  C_56_S_0_L_3_out, I4 =>  C_56_S_0_L_4_out, I5 =>  C_56_S_0_L_5_out); 
C_56_S_1_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_56_S_1_out, I0 =>  C_56_S_1_L_0_out, I1 =>  C_56_S_1_L_1_out, I2 =>  C_56_S_1_L_2_out, I3 =>  C_56_S_1_L_3_out, I4 =>  C_56_S_1_L_4_out, I5 =>  C_56_S_1_L_5_out); 
C_56_S_2_inst : LUT6 generic map(INIT => "1111111011111000111010001110000011111000111010001110000010000000") port map( O =>C_56_S_2_out, I0 =>  C_56_S_2_L_0_out, I1 =>  C_56_S_2_L_1_out, I2 =>  C_56_S_2_L_2_out, I3 =>  C_56_S_2_L_3_out, I4 =>  C_56_S_2_L_4_out, I5 =>  C_56_S_2_L_5_out); 
C_56_S_3_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_56_S_3_out, I0 =>  C_56_S_3_L_0_out, I1 =>  C_56_S_3_L_1_out, I2 =>  C_56_S_3_L_2_out, I3 =>  C_56_S_3_L_3_out, I4 =>  C_56_S_3_L_4_out, I5 =>  C_56_S_3_L_5_out); 
C_56_S_4_inst : LUT6 generic map(INIT => "1111111111111110111111101100100011101100100000001000000000000000") port map( O =>C_56_S_4_out, I0 =>  C_56_S_4_L_0_out, I1 =>  C_56_S_4_L_1_out, I2 =>  C_56_S_4_L_2_out, I3 =>  C_56_S_4_L_3_out, I4 =>  C_56_S_4_L_4_out, I5 =>  C_56_S_4_L_5_out); 
C_56_S_5_inst : LUT6 generic map(INIT => "1111111111111000111111101000000011111110100000001110000000000000") port map( O =>C_56_S_5_out, I0 =>  C_56_S_5_L_0_out, I1 =>  C_56_S_5_L_1_out, I2 =>  C_56_S_5_L_2_out, I3 =>  C_56_S_5_L_3_out, I4 =>  C_56_S_5_L_4_out, I5 =>  C_56_S_5_L_5_out); 

C_56_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_56_out, I0 =>  C_56_S_0_out, I1 =>  C_56_S_1_out, I2 =>  C_56_S_2_out, I3 =>  C_56_S_3_out, I4 =>  C_56_S_4_out, I5 =>  C_56_S_5_out); 

 
C_57_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_57_S_0_out, I0 =>  C_57_S_0_L_0_out, I1 =>  C_57_S_0_L_1_out, I2 =>  C_57_S_0_L_2_out, I3 =>  C_57_S_0_L_3_out, I4 =>  C_57_S_0_L_4_out, I5 =>  C_57_S_0_L_5_out); 
C_57_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010101000000011111110101010001110100010000000") port map( O =>C_57_S_1_out, I0 =>  C_57_S_1_L_0_out, I1 =>  C_57_S_1_L_1_out, I2 =>  C_57_S_1_L_2_out, I3 =>  C_57_S_1_L_3_out, I4 =>  C_57_S_1_L_4_out, I5 =>  C_57_S_1_L_5_out); 
C_57_S_2_inst : LUT6 generic map(INIT => "1111111011111100111111001100100011101100110000001100000010000000") port map( O =>C_57_S_2_out, I0 =>  C_57_S_2_L_0_out, I1 =>  C_57_S_2_L_1_out, I2 =>  C_57_S_2_L_2_out, I3 =>  C_57_S_2_L_3_out, I4 =>  C_57_S_2_L_4_out, I5 =>  C_57_S_2_L_5_out); 
C_57_S_3_inst : LUT6 generic map(INIT => "1111111111111110111111001100000011111100110000001000000000000000") port map( O =>C_57_S_3_out, I0 =>  C_57_S_3_L_0_out, I1 =>  C_57_S_3_L_1_out, I2 =>  C_57_S_3_L_2_out, I3 =>  C_57_S_3_L_3_out, I4 =>  C_57_S_3_L_4_out, I5 =>  C_57_S_3_L_5_out); 
C_57_S_4_inst : LUT6 generic map(INIT => "1111111011111010111010001010000011111010111010001010000010000000") port map( O =>C_57_S_4_out, I0 =>  C_57_S_4_L_0_out, I1 =>  C_57_S_4_L_1_out, I2 =>  C_57_S_4_L_2_out, I3 =>  C_57_S_4_L_3_out, I4 =>  C_57_S_4_L_4_out, I5 =>  C_57_S_4_L_5_out); 
C_57_S_5_inst : LUT6 generic map(INIT => "1111111011101010111010101010100011101010101010001010100010000000") port map( O =>C_57_S_5_out, I0 =>  C_57_S_5_L_0_out, I1 =>  C_57_S_5_L_1_out, I2 =>  C_57_S_5_L_2_out, I3 =>  C_57_S_5_L_3_out, I4 =>  C_57_S_5_L_4_out, I5 =>  C_57_S_5_L_5_out); 

C_57_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_57_out, I0 =>  C_57_S_0_out, I1 =>  C_57_S_1_out, I2 =>  C_57_S_2_out, I3 =>  C_57_S_3_out, I4 =>  C_57_S_4_out, I5 =>  C_57_S_5_out); 

 
C_58_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_58_S_0_out, I0 =>  C_58_S_0_L_0_out, I1 =>  C_58_S_0_L_1_out, I2 =>  C_58_S_0_L_2_out, I3 =>  C_58_S_0_L_3_out, I4 =>  C_58_S_0_L_4_out, I5 =>  C_58_S_0_L_5_out); 
C_58_S_1_inst : LUT6 generic map(INIT => "1110111011101010111010101010100011101010101010001010100010001000") port map( O =>C_58_S_1_out, I0 =>  C_58_S_1_L_0_out, I1 =>  C_58_S_1_L_1_out, I2 =>  C_58_S_1_L_2_out, I3 =>  C_58_S_1_L_3_out, I4 =>  C_58_S_1_L_4_out, I5 =>  C_58_S_1_L_5_out); 
C_58_S_2_inst : LUT6 generic map(INIT => "1111111011111000111111001110000011111000110000001110000010000000") port map( O =>C_58_S_2_out, I0 =>  C_58_S_2_L_0_out, I1 =>  C_58_S_2_L_1_out, I2 =>  C_58_S_2_L_2_out, I3 =>  C_58_S_2_L_3_out, I4 =>  C_58_S_2_L_4_out, I5 =>  C_58_S_2_L_5_out); 
C_58_S_3_inst : LUT6 generic map(INIT => "1111111111101100111111101100000011111100100000001100100000000000") port map( O =>C_58_S_3_out, I0 =>  C_58_S_3_L_0_out, I1 =>  C_58_S_3_L_1_out, I2 =>  C_58_S_3_L_2_out, I3 =>  C_58_S_3_L_3_out, I4 =>  C_58_S_3_L_4_out, I5 =>  C_58_S_3_L_5_out); 
C_58_S_4_inst : LUT6 generic map(INIT => "1111111011111100111110001110100011101000111000001100000010000000") port map( O =>C_58_S_4_out, I0 =>  C_58_S_4_L_0_out, I1 =>  C_58_S_4_L_1_out, I2 =>  C_58_S_4_L_2_out, I3 =>  C_58_S_4_L_3_out, I4 =>  C_58_S_4_L_4_out, I5 =>  C_58_S_4_L_5_out); 
C_58_S_5_inst : LUT6 generic map(INIT => "1111111011101000111011101100100011101100100010001110100010000000") port map( O =>C_58_S_5_out, I0 =>  C_58_S_5_L_0_out, I1 =>  C_58_S_5_L_1_out, I2 =>  C_58_S_5_L_2_out, I3 =>  C_58_S_5_L_3_out, I4 =>  C_58_S_5_L_4_out, I5 =>  C_58_S_5_L_5_out); 

C_58_inst : LUT6 generic map(INIT => "1110101010101010101010101010101010101010101010101010101010101000") port map( O =>C_58_out, I0 =>  C_58_S_0_out, I1 =>  C_58_S_1_out, I2 =>  C_58_S_2_out, I3 =>  C_58_S_3_out, I4 =>  C_58_S_4_out, I5 =>  C_58_S_5_out); 

 
C_59_S_0_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_59_S_0_out, I0 =>  C_59_S_0_L_0_out, I1 =>  C_59_S_0_L_1_out, I2 =>  C_59_S_0_L_2_out, I3 =>  C_59_S_0_L_3_out, I4 =>  C_59_S_0_L_4_out, I5 =>  C_59_S_0_L_5_out); 
C_59_S_1_inst : LUT6 generic map(INIT => "1111111011101000111010001000100011101110111010001110100010000000") port map( O =>C_59_S_1_out, I0 =>  C_59_S_1_L_0_out, I1 =>  C_59_S_1_L_1_out, I2 =>  C_59_S_1_L_2_out, I3 =>  C_59_S_1_L_3_out, I4 =>  C_59_S_1_L_4_out, I5 =>  C_59_S_1_L_5_out); 
C_59_S_2_inst : LUT6 generic map(INIT => "1111111011101000111010001000000011111110111010001110100010000000") port map( O =>C_59_S_2_out, I0 =>  C_59_S_2_L_0_out, I1 =>  C_59_S_2_L_1_out, I2 =>  C_59_S_2_L_2_out, I3 =>  C_59_S_2_L_3_out, I4 =>  C_59_S_2_L_4_out, I5 =>  C_59_S_2_L_5_out); 
C_59_S_3_inst : LUT6 generic map(INIT => "1111111111101010111010101010000011111010101010001010100000000000") port map( O =>C_59_S_3_out, I0 =>  C_59_S_3_L_0_out, I1 =>  C_59_S_3_L_1_out, I2 =>  C_59_S_3_L_2_out, I3 =>  C_59_S_3_L_3_out, I4 =>  C_59_S_3_L_4_out, I5 =>  C_59_S_3_L_5_out); 
C_59_S_4_inst : LUT6 generic map(INIT => "1111111011111000111110001110000011111000111000001110000010000000") port map( O =>C_59_S_4_out, I0 =>  C_59_S_4_L_0_out, I1 =>  C_59_S_4_L_1_out, I2 =>  C_59_S_4_L_2_out, I3 =>  C_59_S_4_L_3_out, I4 =>  C_59_S_4_L_4_out, I5 =>  C_59_S_4_L_5_out); 
C_59_S_5_inst : LUT6 generic map(INIT => "1111111111101110111111101110100011101000100000001000100000000000") port map( O =>C_59_S_5_out, I0 =>  C_59_S_5_L_0_out, I1 =>  C_59_S_5_L_1_out, I2 =>  C_59_S_5_L_2_out, I3 =>  C_59_S_5_L_3_out, I4 =>  C_59_S_5_L_4_out, I5 =>  C_59_S_5_L_5_out); 

C_59_inst : LUT6 generic map(INIT => "1010101010101010101010101010101010101010101010101010101010101010") port map( O =>C_59_out, I0 =>  C_59_S_0_out, I1 =>  C_59_S_1_out, I2 =>  C_59_S_2_out, I3 =>  C_59_S_3_out, I4 =>  C_59_S_4_out, I5 =>  C_59_S_5_out); 

C_0_B_0_inst : LUT6 generic map(INIT => "1001100111001100011001100011001101001110011001111001100111001100") port map( O =>C_0_B_0_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_1_inst : LUT6 generic map(INIT => "1110000111110000100001111100001100001111100001110001111000001111") port map( O =>C_0_B_1_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_2_inst : LUT6 generic map(INIT => "1100001000111100110001000011111101001100001110111101110000110011") port map( O =>C_0_B_2_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_3_inst : LUT6 generic map(INIT => "0101100110011010101000100110011000101010011001100100010110011001") port map( O =>C_0_B_3_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_4_inst : LUT6 generic map(INIT => "0110001000100011110001000100010000110011101110110110011000100010") port map( O =>C_0_B_4_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_5_inst : LUT6 generic map(INIT => "0010100110010110010100100010110100010110011010010010110110010110") port map( O =>C_0_B_5_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_6_inst : LUT6 generic map(INIT => "0001011101111110001111101110110000000001000101110001001101111110") port map( O =>C_0_B_6_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 
C_0_B_7_inst : LUT6 generic map(INIT => "1111111111111110111111101110110011111111111111111111111111111110") port map( O =>C_0_B_7_out, I0 =>  C_0_out, I1 =>  C_1_out, I2 =>  C_2_out, I3 =>  C_3_out, I4 =>  C_4_out, I5 =>  C_5_out); 

C_1_B_0_inst : LUT6 generic map(INIT => "0000000111110000000011111111000010100101000011111111000000001111") port map( O =>C_1_B_0_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_1_inst : LUT6 generic map(INIT => "1010000010100101101010101010010100001010101010100101101010101010") port map( O =>C_1_B_1_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_2_inst : LUT6 generic map(INIT => "1111000011111010000011110000010111110000111100000101111100001111") port map( O =>C_1_B_2_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_3_inst : LUT6 generic map(INIT => "0110000010011001011010011001110010011001011001101100011001101001") port map( O =>C_1_B_3_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_4_inst : LUT6 generic map(INIT => "0001000001111000111010001000001110000111000111100011111011101000") port map( O =>C_1_B_4_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_5_inst : LUT6 generic map(INIT => "0000000011110111111001110111000010001111111100011111000100011000") port map( O =>C_1_B_5_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_6_inst : LUT6 generic map(INIT => "0000000000000000000100001111111101110000111111111111111100001000") port map( O =>C_1_B_6_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 
C_1_B_7_inst : LUT6 generic map(INIT => "1111111111111111111111111111111111111111111111111111111100001000") port map( O =>C_1_B_7_out, I0 =>  C_6_out, I1 =>  C_7_out, I2 =>  C_8_out, I3 =>  C_9_out, I4 =>  C_10_out, I5 =>  C_11_out); 

C_2_B_0_inst : LUT6 generic map(INIT => "1000110011100110000110011001100111000110011001101001100110011000") port map( O =>C_2_B_0_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_1_inst : LUT6 generic map(INIT => "1001100101101110100010000111011110010001111011101000100001110110") port map( O =>C_2_B_1_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_2_inst : LUT6 generic map(INIT => "0100010011011101101110110011001110110011001000100100010011001101") port map( O =>C_2_B_2_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_3_inst : LUT6 generic map(INIT => "1001100101100110001000100101010100101010010001000110011010011001") port map( O =>C_2_B_3_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_4_inst : LUT6 generic map(INIT => "0001000110001000001100111001100111001100011101111000100011101110") port map( O =>C_2_B_4_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_5_inst : LUT6 generic map(INIT => "1101001000111100111100000010110111000011101101001100001100111100") port map( O =>C_2_B_5_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_6_inst : LUT6 generic map(INIT => "1110110011000000110011001100000111111100110010001111110011000000") port map( O =>C_2_B_6_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 
C_2_B_7_inst : LUT6 generic map(INIT => "0000000000000000000000000000000100000000000000000000000000000000") port map( O =>C_2_B_7_out, I0 =>  C_12_out, I1 =>  C_13_out, I2 =>  C_14_out, I3 =>  C_15_out, I4 =>  C_16_out, I5 =>  C_17_out); 

C_3_B_0_inst : LUT6 generic map(INIT => "1000011110100111111110000101100000001110100001111111000101111000") port map( O =>C_3_B_0_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_1_inst : LUT6 generic map(INIT => "1100101111001011101100111001001111000011110010110011001010110011") port map( O =>C_3_B_1_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_2_inst : LUT6 generic map(INIT => "1100000011000000100011110010111111000000110000000000111100001111") port map( O =>C_3_B_2_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_3_inst : LUT6 generic map(INIT => "1101011001010110111010010110100101010110010101100110100101101001") port map( O =>C_3_B_3_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_4_inst : LUT6 generic map(INIT => "1110101110010100110000101011110110010100011010111011110101000010") port map( O =>C_3_B_4_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_5_inst : LUT6 generic map(INIT => "1100111111011011110011111111001000100100010011110000110101001111") port map( O =>C_3_B_5_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_6_inst : LUT6 generic map(INIT => "1111110011101100111111001100110011001000100000111100000110000011") port map( O =>C_3_B_6_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 
C_3_B_7_inst : LUT6 generic map(INIT => "0000000000000000000000000000000000000000000000110000000100000011") port map( O =>C_3_B_7_out, I0 =>  C_18_out, I1 =>  C_19_out, I2 =>  C_20_out, I3 =>  C_21_out, I4 =>  C_22_out, I5 =>  C_23_out); 

C_4_B_0_inst : LUT6 generic map(INIT => "1100111111001111111100000000111100001111000011111111000011110000") port map( O =>C_4_B_0_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_1_inst : LUT6 generic map(INIT => "1111111111111111111100001111111100000000000000000000111100001111") port map( O =>C_4_B_1_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_2_inst : LUT6 generic map(INIT => "1101111011011110010101010101101010100101101001011010010110100101") port map( O =>C_4_B_2_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_3_inst : LUT6 generic map(INIT => "1101111111101100010101011010000011111010000001011111101000000101") port map( O =>C_4_B_3_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_4_inst : LUT6 generic map(INIT => "1110110011111111101010101111111100000000111110100000000011111010") port map( O =>C_4_B_4_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_5_inst : LUT6 generic map(INIT => "1100110011001100000000000000000011111111111111111111111111111111") port map( O =>C_4_B_5_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_6_inst : LUT6 generic map(INIT => "1111111111111111110011001100110011001100110011000011001100110011") port map( O =>C_4_B_6_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 
C_4_B_7_inst : LUT6 generic map(INIT => "0000000000000000000000000000000000000000000000000011001100110011") port map( O =>C_4_B_7_out, I0 =>  C_24_out, I1 =>  C_25_out, I2 =>  C_26_out, I3 =>  C_27_out, I4 =>  C_28_out, I5 =>  C_29_out); 

C_5_B_0_inst : LUT6 generic map(INIT => "1001111000001111111110001001111011110000110110101110000111110000") port map( O =>C_5_B_0_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_1_inst : LUT6 generic map(INIT => "1001011110010110100100011001011111100110111011001111011011100110") port map( O =>C_5_B_1_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_2_inst : LUT6 generic map(INIT => "1000000101111110111110001000000110011110111010011110000110011110") port map( O =>C_5_B_2_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_3_inst : LUT6 generic map(INIT => "1100001111000010101110111100001111000010110101001010001111000010") port map( O =>C_5_B_3_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_4_inst : LUT6 generic map(INIT => "1000110011110010110010111000110011110010100011111010110011110010") port map( O =>C_5_B_4_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_5_inst : LUT6 generic map(INIT => "1011001111000001101101111011001110111110101100111110110010111110") port map( O =>C_5_B_5_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_6_inst : LUT6 generic map(INIT => "1110100110101001111010011110100111101000111010011111101011101000") port map( O =>C_5_B_6_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 
C_5_B_7_inst : LUT6 generic map(INIT => "0000000100000001000000010000000100000000000000010000000000000000") port map( O =>C_5_B_7_out, I0 =>  C_30_out, I1 =>  C_31_out, I2 =>  C_32_out, I3 =>  C_33_out, I4 =>  C_34_out, I5 =>  C_35_out); 

C_6_B_0_inst : LUT6 generic map(INIT => "1011010011010110011010011001010001000010011010011001011001001011") port map( O =>C_6_B_0_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_1_inst : LUT6 generic map(INIT => "1100100000010111100000010001011110000011011111100001011101111100") port map( O =>C_6_B_1_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_2_inst : LUT6 generic map(INIT => "1100110011011011001100100010010011001111101100110010010001001100") port map( O =>C_6_B_2_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_3_inst : LUT6 generic map(INIT => "1111000000011100001111001100011111110011001111000011100010001111") port map( O =>C_6_B_3_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_4_inst : LUT6 generic map(INIT => "1001100101111001010110010110000101100101101001101010011010010110") port map( O =>C_6_B_4_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_5_inst : LUT6 generic map(INIT => "1101110101011101010111010100010110111010111110111111101111011011") port map( O =>C_6_B_5_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_6_inst : LUT6 generic map(INIT => "0100010011000100110001001101110010011001100110011001100110111001") port map( O =>C_6_B_6_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 
C_6_B_7_inst : LUT6 generic map(INIT => "1111111111111111111111111111111110111011101110111011101110111011") port map( O =>C_6_B_7_out, I0 =>  C_36_out, I1 =>  C_37_out, I2 =>  C_38_out, I3 =>  C_39_out, I4 =>  C_40_out, I5 =>  C_41_out); 

C_7_B_0_inst : LUT6 generic map(INIT => "1100110100110011111111110010001011001101001100111111111100100000") port map( O =>C_7_B_0_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_1_inst : LUT6 generic map(INIT => "0011110011110000110000110001111000111100111100001100001100011100") port map( O =>C_7_B_1_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_2_inst : LUT6 generic map(INIT => "0011000011000011111100111100110100110000110000111111001111001111") port map( O =>C_7_B_2_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_3_inst : LUT6 generic map(INIT => "1100111100001100000011000000000011001111000011000000110000000000") port map( O =>C_7_B_3_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_4_inst : LUT6 generic map(INIT => "0011001100110011001100110011001100110011001100110011001100110011") port map( O =>C_7_B_4_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_5_inst : LUT6 generic map(INIT => "1111111100000000000000001111111111111111000000000000000011111111") port map( O =>C_7_B_5_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_6_inst : LUT6 generic map(INIT => "0000000000000000111111110000000011111111111111110000000011111111") port map( O =>C_7_B_6_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 
C_7_B_7_inst : LUT6 generic map(INIT => "0000000000000000000000000000000011111111111111110000000011111111") port map( O =>C_7_B_7_out, I0 =>  C_42_out, I1 =>  C_43_out, I2 =>  C_44_out, I3 =>  C_45_out, I4 =>  C_46_out, I5 =>  C_47_out); 

C_8_B_0_inst : LUT6 generic map(INIT => "1000111101110000111100010000111000001100111000111110011100111000") port map( O =>C_8_B_0_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_1_inst : LUT6 generic map(INIT => "1011001100111100001111001100110100110000001011000010110011001011") port map( O =>C_8_B_1_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_2_inst : LUT6 generic map(INIT => "0100001111000000001111110000111111000000110100000010111100001011") port map( O =>C_8_B_2_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_3_inst : LUT6 generic map(INIT => "1001010110010110101010011001100110010110100101101011100110011101") port map( O =>C_8_B_3_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_4_inst : LUT6 generic map(INIT => "0010101011010100000000101101110111010100001010111111110100100010") port map( O =>C_8_B_4_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_5_inst : LUT6 generic map(INIT => "1001011010111101100101101011010010111101011010011001010001101001") port map( O =>C_8_B_5_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_6_inst : LUT6 generic map(INIT => "1101010011010110110101001101011000101001101111010010100110111101") port map( O =>C_8_B_6_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 
C_8_B_7_inst : LUT6 generic map(INIT => "1101010011010100110101001101010011111101111111011111110111111101") port map( O =>C_8_B_7_out, I0 =>  C_48_out, I1 =>  C_49_out, I2 =>  C_50_out, I3 =>  C_51_out, I4 =>  C_52_out, I5 =>  C_53_out); 

C_9_B_0_inst : LUT6 generic map(INIT => "0001000011110111000000000111011110101010000100011010111000010000") port map( O =>C_9_B_0_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_1_inst : LUT6 generic map(INIT => "1000011001100001100101001110000101101001011110000110100101111001") port map( O =>C_9_B_1_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_2_inst : LUT6 generic map(INIT => "1000111000010000011100011110111111100111000010000001100011110111") port map( O =>C_9_B_2_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_3_inst : LUT6 generic map(INIT => "1110011101101001100101001000011010000110011000011001111010010110") port map( O =>C_9_B_3_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_4_inst : LUT6 generic map(INIT => "0110000100011000100011000110000110011110111001110111100110001110") port map( O =>C_9_B_4_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_5_inst : LUT6 generic map(INIT => "1101110011000100010000000010001101000010001000110011101110111101") port map( O =>C_9_B_5_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_6_inst : LUT6 generic map(INIT => "0000000011111111000000001101110011111101001000111100010010111111") port map( O =>C_9_B_6_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 
C_9_B_7_inst : LUT6 generic map(INIT => "1111111111111111111111111111111111111111001000111111111110111111") port map( O =>C_9_B_7_out, I0 =>  C_54_out, I1 =>  C_55_out, I2 =>  C_56_out, I3 =>  C_57_out, I4 =>  C_58_out, I5 =>  C_59_out); 


out_fin <= C_0_B_7_out  & C_0_B_6_out  & C_0_B_5_out  & C_0_B_4_out  & C_0_B_3_out  & C_0_B_2_out  & C_0_B_1_out  & C_0_B_0_out  & C_1_B_7_out  & C_1_B_6_out  & C_1_B_5_out  & C_1_B_4_out  & C_1_B_3_out  & C_1_B_2_out  & C_1_B_1_out  & C_1_B_0_out  & C_2_B_7_out  & C_2_B_6_out  & C_2_B_5_out  & C_2_B_4_out  & C_2_B_3_out  & C_2_B_2_out  & C_2_B_1_out  & C_2_B_0_out  & C_3_B_7_out  & C_3_B_6_out  & C_3_B_5_out  & C_3_B_4_out  & C_3_B_3_out  & C_3_B_2_out  & C_3_B_1_out  & C_3_B_0_out  & C_4_B_7_out  & C_4_B_6_out  & C_4_B_5_out  & C_4_B_4_out  & C_4_B_3_out  & C_4_B_2_out  & C_4_B_1_out  & C_4_B_0_out  & C_5_B_7_out  & C_5_B_6_out  & C_5_B_5_out  & C_5_B_4_out  & C_5_B_3_out  & C_5_B_2_out  & C_5_B_1_out  & C_5_B_0_out  & C_6_B_7_out  & C_6_B_6_out  & C_6_B_5_out  & C_6_B_4_out  & C_6_B_3_out  & C_6_B_2_out  & C_6_B_1_out  & C_6_B_0_out  & C_7_B_7_out  & C_7_B_6_out  & C_7_B_5_out  & C_7_B_4_out  & C_7_B_3_out  & C_7_B_2_out  & C_7_B_1_out  & C_7_B_0_out  & C_8_B_7_out  & C_8_B_6_out  & C_8_B_5_out  & C_8_B_4_out  & C_8_B_3_out  & C_8_B_2_out  & C_8_B_1_out  & C_8_B_0_out  & C_9_B_7_out  & C_9_B_6_out  & C_9_B_5_out  & C_9_B_4_out  & C_9_B_3_out  & C_9_B_2_out  & C_9_B_1_out  & C_9_B_0_out ; 
--cor_out <= cor_in;
--pred_out <= C_0_out &C_1_out &C_2_out &C_3_out &C_4_out &C_5_out &C_6_out &C_7_out &C_8_out &C_9_out &C_10_out &C_11_out &C_12_out &C_13_out &C_14_out &C_15_out &C_16_out &C_17_out &C_18_out &C_19_out &C_20_out &C_21_out &C_22_out &C_23_out &C_24_out &C_25_out &C_26_out &C_27_out &C_28_out &C_29_out &C_30_out &C_31_out &C_32_out &C_33_out &C_34_out &C_35_out &C_36_out &C_37_out &C_38_out &C_39_out &C_40_out &C_41_out &C_42_out &C_43_out &C_44_out &C_45_out &C_46_out &C_47_out &C_48_out &C_49_out &C_50_out &C_51_out &C_52_out &C_53_out &C_54_out &C_55_out &C_56_out &C_57_out &C_58_out &C_59_out ; 

end Behavioral;

