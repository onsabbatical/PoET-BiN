--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:20:18 07/23/2019
-- Design Name:   
-- Module Name:   D:/siva/Masters/Thesis/07_ETE_19/part_svhn/cifar_fin_layer_tb.vhd
-- Project Name:  part_svhn
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: cifar_fin_layer
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY cifar_fin_layer_tb IS
END cifar_fin_layer_tb;
 
ARCHITECTURE behavior OF cifar_fin_layer_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT cifar_fin_layer
    PORT(
         inp_feat : IN  std_logic_vector(79 downto 0);
         cor_in : IN  std_logic_vector(79 downto 0);
         cor_out : OUT  std_logic_vector(79 downto 0);
         out_fin : OUT  std_logic_vector(79 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal inp_feat : std_logic_vector(79 downto 0) := (others => '0');
   signal cor_in : std_logic_vector(79 downto 0) := (others => '0');

 	--Outputs
   signal cor_out : std_logic_vector(79 downto 0);
   signal out_fin : std_logic_vector(79 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: cifar_fin_layer PORT MAP (
          inp_feat => inp_feat,
          cor_in => cor_in,
          cor_out => cor_out,
          out_fin => out_fin
        );

   -- Clock process definitions
   --<clock>_process :process
   --begin
	--	<clock> <= '0';
	--	wait for <clock>_period/2;
	--	<clock> <= '1';
	--	wait for <clock>_period/2;
   -- end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

     -- wait for <clock>_period*10;
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010101000000011";cor_in <= "11011111110101111110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010101010100011";cor_in <= "11100001110101111110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111011101000100000011";cor_in <= "11011111001000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111011101000100000011";cor_in <= "11011111001000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111011010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111010111011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111011010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000100011";cor_in <= "11010100111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101010101010010100010110010000101011111010010111000111011";cor_in <= "11010010111000001110000011011111111000001101111111010000001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010101101001110000101011111010010111010000100";cor_in <= "00011010111000001110000011011111001000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010101101001110000101011111010010111000000011";cor_in <= "11011111111000001110000011011111001000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101111001011101001110000101011111010010111000000011";cor_in <= "11011111111000001110000011011111001000000001000111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010101101001110000101011111010010111000000011";cor_in <= "11011111111000001110000011011111001000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111011101000100000011";cor_in <= "11011111001000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101011010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010101101001110000101011111010010111000000011";cor_in <= "11011111111000001110000011011111001000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "00010010101110000100011001010101010010100010110010000101011111011100000100010010";cor_in <= "11101000000110111110000011011111111000001101111111010000110111101110000000000000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111011010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101100010010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000000000011011010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011001010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111100010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101010101011010100010110010000100011111010010111000000011";cor_in <= "11011111111000001110000011010110111000001101111111010000001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110011000101011111010010111000000011";cor_in <= "11011111111000001110000011100110111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110011000101011111010010111000000011";cor_in <= "11011111111000001110000011100110111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111011010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101011010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111011101000100000011";cor_in <= "11011111001000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111011010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010100101001011010010111000000011";cor_in <= "11011111111000001111011011101001111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111011101000100000011";cor_in <= "11011111001000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111011101000100000011";cor_in <= "11011111001000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101101101010010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000000001111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101100000100010111000000011";cor_in <= "11011111111000000010000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110011001100011111010010111000110011";cor_in <= "11001101111000001110000011011101111000001101111111011010001000001110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "10000011101110000100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111101110000000100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001011101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111011010110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110001111010011111010010111000000011";cor_in <= "11011111111000001110000000011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100010001110100011001010101010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111111010000110111100011101111100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010101101001110000101011111010010111000000011";cor_in <= "11011111111000001110000011011111001000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011010101010010010100010110010000101011111010010111000000011";cor_in <= "11011111111000001110000011011111111000001101111100100000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110000100011001010101010010100010110010000101011111010010111011111100";cor_in <= "00100000111000001110000011011111111000001101111111010000110111101110000011100000" ; wait for 10 ns; 
inp_feat <= "01111100101110001011100101011101010010100010110010000101011111010010111000011011";cor_in <= "11011101111000001110000011011111111000001101111111011010001000001110000011100000" ; wait for 10 ns; 

      -- insert stimulus here 

      wait;
   end process;

END;
